// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 15.1.0 Build 185 10/21/2015 SJ Lite Edition"

// DATE "07/21/2017 00:34:00"

// 
// Device: Altera 5CSEMA5F31C6 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module sine (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	clk,
	clken,
	phi_inc_i,
	freq_mod_i,
	phase_mod_i,
	fsin_o,
	out_valid,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	clk;
input 	clken;
input 	[31:0] phi_inc_i;
input 	[31:0] freq_mod_i;
input 	[15:0] phase_mod_i;
output 	[23:0] fsin_o;
output 	out_valid;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \nco_ii_0|ux710isdr|data_ready~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[20]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[21]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[22]~q ;
wire \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[23]~q ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \clk~input_o ;
wire \clken~input_o ;
wire \reset_n~input_o ;
wire \phase_mod_i[8]~input_o ;
wire \phase_mod_i[9]~input_o ;
wire \phase_mod_i[10]~input_o ;
wire \phase_mod_i[11]~input_o ;
wire \phase_mod_i[12]~input_o ;
wire \phase_mod_i[13]~input_o ;
wire \phase_mod_i[14]~input_o ;
wire \phase_mod_i[15]~input_o ;
wire \phase_mod_i[0]~input_o ;
wire \phase_mod_i[1]~input_o ;
wire \phase_mod_i[2]~input_o ;
wire \phase_mod_i[3]~input_o ;
wire \phase_mod_i[4]~input_o ;
wire \phase_mod_i[5]~input_o ;
wire \phase_mod_i[6]~input_o ;
wire \phase_mod_i[7]~input_o ;
wire \freq_mod_i[24]~input_o ;
wire \phi_inc_i[24]~input_o ;
wire \freq_mod_i[25]~input_o ;
wire \phi_inc_i[25]~input_o ;
wire \freq_mod_i[26]~input_o ;
wire \phi_inc_i[26]~input_o ;
wire \freq_mod_i[27]~input_o ;
wire \phi_inc_i[27]~input_o ;
wire \freq_mod_i[28]~input_o ;
wire \phi_inc_i[28]~input_o ;
wire \freq_mod_i[29]~input_o ;
wire \phi_inc_i[29]~input_o ;
wire \freq_mod_i[30]~input_o ;
wire \phi_inc_i[30]~input_o ;
wire \freq_mod_i[31]~input_o ;
wire \phi_inc_i[31]~input_o ;
wire \freq_mod_i[16]~input_o ;
wire \phi_inc_i[16]~input_o ;
wire \freq_mod_i[17]~input_o ;
wire \phi_inc_i[17]~input_o ;
wire \freq_mod_i[18]~input_o ;
wire \phi_inc_i[18]~input_o ;
wire \freq_mod_i[19]~input_o ;
wire \phi_inc_i[19]~input_o ;
wire \freq_mod_i[20]~input_o ;
wire \phi_inc_i[20]~input_o ;
wire \freq_mod_i[21]~input_o ;
wire \phi_inc_i[21]~input_o ;
wire \freq_mod_i[22]~input_o ;
wire \phi_inc_i[22]~input_o ;
wire \freq_mod_i[23]~input_o ;
wire \phi_inc_i[23]~input_o ;
wire \freq_mod_i[15]~input_o ;
wire \phi_inc_i[15]~input_o ;
wire \freq_mod_i[14]~input_o ;
wire \phi_inc_i[14]~input_o ;
wire \freq_mod_i[13]~input_o ;
wire \phi_inc_i[13]~input_o ;
wire \freq_mod_i[12]~input_o ;
wire \phi_inc_i[12]~input_o ;
wire \freq_mod_i[11]~input_o ;
wire \phi_inc_i[11]~input_o ;
wire \freq_mod_i[10]~input_o ;
wire \phi_inc_i[10]~input_o ;
wire \freq_mod_i[9]~input_o ;
wire \phi_inc_i[9]~input_o ;
wire \freq_mod_i[8]~input_o ;
wire \phi_inc_i[8]~input_o ;
wire \freq_mod_i[7]~input_o ;
wire \phi_inc_i[7]~input_o ;
wire \freq_mod_i[6]~input_o ;
wire \phi_inc_i[6]~input_o ;
wire \freq_mod_i[5]~input_o ;
wire \phi_inc_i[5]~input_o ;
wire \freq_mod_i[4]~input_o ;
wire \phi_inc_i[4]~input_o ;
wire \freq_mod_i[3]~input_o ;
wire \phi_inc_i[3]~input_o ;
wire \freq_mod_i[2]~input_o ;
wire \phi_inc_i[2]~input_o ;
wire \freq_mod_i[1]~input_o ;
wire \phi_inc_i[1]~input_o ;
wire \freq_mod_i[0]~input_o ;
wire \phi_inc_i[0]~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TDIUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ;
wire \nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|Equal2~2_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ;
wire \nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ;
wire \nabboc|pzdyqx_impl_inst|AMGP4450~q ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0_combout ;
wire \nabboc|pzdyqx_impl_inst|comb~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ;
wire \nabboc|pzdyqx_impl_inst|sdr~combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ;
wire \nabboc|pzdyqx_impl_inst|dr_scan~combout ;
wire \nabboc|pzdyqx_impl_inst|KNOR6738~q ;
wire \nabboc|pzdyqx_impl_inst|tdo~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;


sine_sine_nco_ii_0 nco_ii_0(
	.data_ready(\nco_ii_0|ux710isdr|data_ready~q ),
	.pipeline_dffe_0(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_15(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_16(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_19(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_20(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_21(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_22(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_23(\nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[23]~q ),
	.GND_port(\~GND~combout ),
	.NJQG9082(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.clk(\clk~input_o ),
	.clken(\clken~input_o ),
	.reset_n(\reset_n~input_o ),
	.phase_mod_i_8(\phase_mod_i[8]~input_o ),
	.phase_mod_i_9(\phase_mod_i[9]~input_o ),
	.phase_mod_i_10(\phase_mod_i[10]~input_o ),
	.phase_mod_i_11(\phase_mod_i[11]~input_o ),
	.phase_mod_i_12(\phase_mod_i[12]~input_o ),
	.phase_mod_i_13(\phase_mod_i[13]~input_o ),
	.phase_mod_i_14(\phase_mod_i[14]~input_o ),
	.phase_mod_i_15(\phase_mod_i[15]~input_o ),
	.phase_mod_i_0(\phase_mod_i[0]~input_o ),
	.phase_mod_i_1(\phase_mod_i[1]~input_o ),
	.phase_mod_i_2(\phase_mod_i[2]~input_o ),
	.phase_mod_i_3(\phase_mod_i[3]~input_o ),
	.phase_mod_i_4(\phase_mod_i[4]~input_o ),
	.phase_mod_i_5(\phase_mod_i[5]~input_o ),
	.phase_mod_i_6(\phase_mod_i[6]~input_o ),
	.phase_mod_i_7(\phase_mod_i[7]~input_o ),
	.freq_mod_i_24(\freq_mod_i[24]~input_o ),
	.phi_inc_i_24(\phi_inc_i[24]~input_o ),
	.freq_mod_i_25(\freq_mod_i[25]~input_o ),
	.phi_inc_i_25(\phi_inc_i[25]~input_o ),
	.freq_mod_i_26(\freq_mod_i[26]~input_o ),
	.phi_inc_i_26(\phi_inc_i[26]~input_o ),
	.freq_mod_i_27(\freq_mod_i[27]~input_o ),
	.phi_inc_i_27(\phi_inc_i[27]~input_o ),
	.freq_mod_i_28(\freq_mod_i[28]~input_o ),
	.phi_inc_i_28(\phi_inc_i[28]~input_o ),
	.freq_mod_i_29(\freq_mod_i[29]~input_o ),
	.phi_inc_i_29(\phi_inc_i[29]~input_o ),
	.freq_mod_i_30(\freq_mod_i[30]~input_o ),
	.phi_inc_i_30(\phi_inc_i[30]~input_o ),
	.freq_mod_i_31(\freq_mod_i[31]~input_o ),
	.phi_inc_i_31(\phi_inc_i[31]~input_o ),
	.freq_mod_i_16(\freq_mod_i[16]~input_o ),
	.phi_inc_i_16(\phi_inc_i[16]~input_o ),
	.freq_mod_i_17(\freq_mod_i[17]~input_o ),
	.phi_inc_i_17(\phi_inc_i[17]~input_o ),
	.freq_mod_i_18(\freq_mod_i[18]~input_o ),
	.phi_inc_i_18(\phi_inc_i[18]~input_o ),
	.freq_mod_i_19(\freq_mod_i[19]~input_o ),
	.phi_inc_i_19(\phi_inc_i[19]~input_o ),
	.freq_mod_i_20(\freq_mod_i[20]~input_o ),
	.phi_inc_i_20(\phi_inc_i[20]~input_o ),
	.freq_mod_i_21(\freq_mod_i[21]~input_o ),
	.phi_inc_i_21(\phi_inc_i[21]~input_o ),
	.freq_mod_i_22(\freq_mod_i[22]~input_o ),
	.phi_inc_i_22(\phi_inc_i[22]~input_o ),
	.freq_mod_i_23(\freq_mod_i[23]~input_o ),
	.phi_inc_i_23(\phi_inc_i[23]~input_o ),
	.freq_mod_i_15(\freq_mod_i[15]~input_o ),
	.phi_inc_i_15(\phi_inc_i[15]~input_o ),
	.freq_mod_i_14(\freq_mod_i[14]~input_o ),
	.phi_inc_i_14(\phi_inc_i[14]~input_o ),
	.freq_mod_i_13(\freq_mod_i[13]~input_o ),
	.phi_inc_i_13(\phi_inc_i[13]~input_o ),
	.freq_mod_i_12(\freq_mod_i[12]~input_o ),
	.phi_inc_i_12(\phi_inc_i[12]~input_o ),
	.freq_mod_i_11(\freq_mod_i[11]~input_o ),
	.phi_inc_i_11(\phi_inc_i[11]~input_o ),
	.freq_mod_i_10(\freq_mod_i[10]~input_o ),
	.phi_inc_i_10(\phi_inc_i[10]~input_o ),
	.freq_mod_i_9(\freq_mod_i[9]~input_o ),
	.phi_inc_i_9(\phi_inc_i[9]~input_o ),
	.freq_mod_i_8(\freq_mod_i[8]~input_o ),
	.phi_inc_i_8(\phi_inc_i[8]~input_o ),
	.freq_mod_i_7(\freq_mod_i[7]~input_o ),
	.phi_inc_i_7(\phi_inc_i[7]~input_o ),
	.freq_mod_i_6(\freq_mod_i[6]~input_o ),
	.phi_inc_i_6(\phi_inc_i[6]~input_o ),
	.freq_mod_i_5(\freq_mod_i[5]~input_o ),
	.phi_inc_i_5(\phi_inc_i[5]~input_o ),
	.freq_mod_i_4(\freq_mod_i[4]~input_o ),
	.phi_inc_i_4(\phi_inc_i[4]~input_o ),
	.freq_mod_i_3(\freq_mod_i[3]~input_o ),
	.phi_inc_i_3(\phi_inc_i[3]~input_o ),
	.freq_mod_i_2(\freq_mod_i[2]~input_o ),
	.phi_inc_i_2(\phi_inc_i[2]~input_o ),
	.freq_mod_i_1(\freq_mod_i[1]~input_o ),
	.phi_inc_i_1(\phi_inc_i[1]~input_o ),
	.freq_mod_i_0(\freq_mod_i[0]~input_o ),
	.phi_inc_i_0(\phi_inc_i[0]~input_o ));

assign \clk~input_o  = clk;

assign \clken~input_o  = clken;

assign \reset_n~input_o  = reset_n;

assign \phase_mod_i[8]~input_o  = phase_mod_i[8];

assign \phase_mod_i[9]~input_o  = phase_mod_i[9];

assign \phase_mod_i[10]~input_o  = phase_mod_i[10];

assign \phase_mod_i[11]~input_o  = phase_mod_i[11];

assign \phase_mod_i[12]~input_o  = phase_mod_i[12];

assign \phase_mod_i[13]~input_o  = phase_mod_i[13];

assign \phase_mod_i[14]~input_o  = phase_mod_i[14];

assign \phase_mod_i[15]~input_o  = phase_mod_i[15];

assign \phase_mod_i[0]~input_o  = phase_mod_i[0];

assign \phase_mod_i[1]~input_o  = phase_mod_i[1];

assign \phase_mod_i[2]~input_o  = phase_mod_i[2];

assign \phase_mod_i[3]~input_o  = phase_mod_i[3];

assign \phase_mod_i[4]~input_o  = phase_mod_i[4];

assign \phase_mod_i[5]~input_o  = phase_mod_i[5];

assign \phase_mod_i[6]~input_o  = phase_mod_i[6];

assign \phase_mod_i[7]~input_o  = phase_mod_i[7];

assign \freq_mod_i[24]~input_o  = freq_mod_i[24];

assign \phi_inc_i[24]~input_o  = phi_inc_i[24];

assign \freq_mod_i[25]~input_o  = freq_mod_i[25];

assign \phi_inc_i[25]~input_o  = phi_inc_i[25];

assign \freq_mod_i[26]~input_o  = freq_mod_i[26];

assign \phi_inc_i[26]~input_o  = phi_inc_i[26];

assign \freq_mod_i[27]~input_o  = freq_mod_i[27];

assign \phi_inc_i[27]~input_o  = phi_inc_i[27];

assign \freq_mod_i[28]~input_o  = freq_mod_i[28];

assign \phi_inc_i[28]~input_o  = phi_inc_i[28];

assign \freq_mod_i[29]~input_o  = freq_mod_i[29];

assign \phi_inc_i[29]~input_o  = phi_inc_i[29];

assign \freq_mod_i[30]~input_o  = freq_mod_i[30];

assign \phi_inc_i[30]~input_o  = phi_inc_i[30];

assign \freq_mod_i[31]~input_o  = freq_mod_i[31];

assign \phi_inc_i[31]~input_o  = phi_inc_i[31];

assign \freq_mod_i[16]~input_o  = freq_mod_i[16];

assign \phi_inc_i[16]~input_o  = phi_inc_i[16];

assign \freq_mod_i[17]~input_o  = freq_mod_i[17];

assign \phi_inc_i[17]~input_o  = phi_inc_i[17];

assign \freq_mod_i[18]~input_o  = freq_mod_i[18];

assign \phi_inc_i[18]~input_o  = phi_inc_i[18];

assign \freq_mod_i[19]~input_o  = freq_mod_i[19];

assign \phi_inc_i[19]~input_o  = phi_inc_i[19];

assign \freq_mod_i[20]~input_o  = freq_mod_i[20];

assign \phi_inc_i[20]~input_o  = phi_inc_i[20];

assign \freq_mod_i[21]~input_o  = freq_mod_i[21];

assign \phi_inc_i[21]~input_o  = phi_inc_i[21];

assign \freq_mod_i[22]~input_o  = freq_mod_i[22];

assign \phi_inc_i[22]~input_o  = phi_inc_i[22];

assign \freq_mod_i[23]~input_o  = freq_mod_i[23];

assign \phi_inc_i[23]~input_o  = phi_inc_i[23];

assign \freq_mod_i[15]~input_o  = freq_mod_i[15];

assign \phi_inc_i[15]~input_o  = phi_inc_i[15];

assign \freq_mod_i[14]~input_o  = freq_mod_i[14];

assign \phi_inc_i[14]~input_o  = phi_inc_i[14];

assign \freq_mod_i[13]~input_o  = freq_mod_i[13];

assign \phi_inc_i[13]~input_o  = phi_inc_i[13];

assign \freq_mod_i[12]~input_o  = freq_mod_i[12];

assign \phi_inc_i[12]~input_o  = phi_inc_i[12];

assign \freq_mod_i[11]~input_o  = freq_mod_i[11];

assign \phi_inc_i[11]~input_o  = phi_inc_i[11];

assign \freq_mod_i[10]~input_o  = freq_mod_i[10];

assign \phi_inc_i[10]~input_o  = phi_inc_i[10];

assign \freq_mod_i[9]~input_o  = freq_mod_i[9];

assign \phi_inc_i[9]~input_o  = phi_inc_i[9];

assign \freq_mod_i[8]~input_o  = freq_mod_i[8];

assign \phi_inc_i[8]~input_o  = phi_inc_i[8];

assign \freq_mod_i[7]~input_o  = freq_mod_i[7];

assign \phi_inc_i[7]~input_o  = phi_inc_i[7];

assign \freq_mod_i[6]~input_o  = freq_mod_i[6];

assign \phi_inc_i[6]~input_o  = phi_inc_i[6];

assign \freq_mod_i[5]~input_o  = freq_mod_i[5];

assign \phi_inc_i[5]~input_o  = phi_inc_i[5];

assign \freq_mod_i[4]~input_o  = freq_mod_i[4];

assign \phi_inc_i[4]~input_o  = phi_inc_i[4];

assign \freq_mod_i[3]~input_o  = freq_mod_i[3];

assign \phi_inc_i[3]~input_o  = phi_inc_i[3];

assign \freq_mod_i[2]~input_o  = freq_mod_i[2];

assign \phi_inc_i[2]~input_o  = phi_inc_i[2];

assign \freq_mod_i[1]~input_o  = freq_mod_i[1];

assign \phi_inc_i[1]~input_o  = phi_inc_i[1];

assign \freq_mod_i[0]~input_o  = freq_mod_i[0];

assign \phi_inc_i[0]~input_o  = phi_inc_i[0];

assign fsin_o[0] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ;

assign fsin_o[1] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ;

assign fsin_o[2] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;

assign fsin_o[3] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;

assign fsin_o[4] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;

assign fsin_o[5] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;

assign fsin_o[6] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;

assign fsin_o[7] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;

assign fsin_o[8] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;

assign fsin_o[9] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;

assign fsin_o[10] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;

assign fsin_o[11] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;

assign fsin_o[12] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;

assign fsin_o[13] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;

assign fsin_o[14] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;

assign fsin_o[15] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;

assign fsin_o[16] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[16]~q ;

assign fsin_o[17] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[17]~q ;

assign fsin_o[18] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[18]~q ;

assign fsin_o[19] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[19]~q ;

assign fsin_o[20] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[20]~q ;

assign fsin_o[21] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[21]~q ;

assign fsin_o[22] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[22]~q ;

assign fsin_o[23] = \nco_ii_0|blk0|lpm_add_sub_component|auto_generated|pipeline_dffe[23]~q ;

assign out_valid = \nco_ii_0|ux710isdr|data_ready~q ;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cyclonev_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 64'h6666666666666666;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 64'h9696969696969696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\~GND~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3 .lut_mask = 64'hF9F6FFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 .lut_mask = 64'hFF96FFFFFF96FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .lut_mask = 64'h7FFFDFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .lut_mask = 64'h6666666666666666;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .lut_mask = 64'h6666666666666666;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .lut_mask = 64'hDEDEDEDEDEDEDEDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .lut_mask = 64'hEDDEEDDEEDDEEDDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .lut_mask = 64'hDEEDEDDEDEEDEDDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .lut_mask = 64'hEDDEDEEDDEEDEDDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .lut_mask = 64'hBEBEBEBEBEBEBEBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .lut_mask = 64'hBEEBEBBEBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .lut_mask = 64'hBEEBEBBEBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|SQHZ7915_1 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_1 .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|SQHZ7915_2 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_2 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 64'hFDF7FFFFF7FDFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 64'hDFD5FFFFDFD5FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|AMGP4450~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|AMGP4450 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|AMGP4450 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|AMGP4450 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|NJQG9082~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|NJQG9082 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 64'hCF5FFFFFCF5FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .lut_mask = 64'hAFFAAFFAAFFAAFFA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .lut_mask = 64'hBEEBBEEBEBBEEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .lut_mask = 64'hFFFFFFBFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 64'hFFFFFFF6FFFFFFF6;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 64'hD1FFD1FFD1FFD1FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .lut_mask = 64'hF7D5F7D5F7D5F7D5;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .lut_mask = 64'hD8FFFFFFD8FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 64'hEFFFFEFFEFFFFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 .lut_mask = 64'hFFEFFFFFFFEFFFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 .lut_mask = 64'hBFEFFFFFBFEFFFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 .lut_mask = 64'hFBFEEBBEFBFEEBBE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|comb~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|comb~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|comb~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \nabboc|pzdyqx_impl_inst|comb~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .lut_mask = 64'h6996F9F66996F9F6;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .lut_mask = 64'hDDF5DFFDDDF5DFFD;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 .lut_mask = 64'h6996F9F66996F9F6;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datae(!\altera_internal_jtag~TDIUTAP ),
	.dataf(!\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 .lut_mask = 64'hB1FFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|sdr (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|sdr .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|sdr .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \nabboc|pzdyqx_impl_inst|sdr .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|dr_scan (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|dr_scan .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|dr_scan .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \nabboc|pzdyqx_impl_inst|dr_scan .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|KNOR6738 (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|tdo~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .lut_mask = 64'hF5F5F5F5F5F5F5F5;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(gnd),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .lut_mask = 64'h5F5FF5F55F5FF5F5;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(gnd),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .lut_mask = 64'hD7D77D7DD7D77D7D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(gnd),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .lut_mask = 64'h7D7DD7D7D7D77D7D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .lut_mask = 64'hD77D7DD77DD7D77D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|~GND .extended_lut = "off";
defparam \auto_hub|~GND .lut_mask = 64'h0000000000000000;
defparam \auto_hub|~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .shared_arith = "off";

endmodule

module sine_sine_nco_ii_0 (
	data_ready,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	GND_port,
	NJQG9082,
	clk,
	clken,
	reset_n,
	phase_mod_i_8,
	phase_mod_i_9,
	phase_mod_i_10,
	phase_mod_i_11,
	phase_mod_i_12,
	phase_mod_i_13,
	phase_mod_i_14,
	phase_mod_i_15,
	phase_mod_i_0,
	phase_mod_i_1,
	phase_mod_i_2,
	phase_mod_i_3,
	phase_mod_i_4,
	phase_mod_i_5,
	phase_mod_i_6,
	phase_mod_i_7,
	freq_mod_i_24,
	phi_inc_i_24,
	freq_mod_i_25,
	phi_inc_i_25,
	freq_mod_i_26,
	phi_inc_i_26,
	freq_mod_i_27,
	phi_inc_i_27,
	freq_mod_i_28,
	phi_inc_i_28,
	freq_mod_i_29,
	phi_inc_i_29,
	freq_mod_i_30,
	phi_inc_i_30,
	freq_mod_i_31,
	phi_inc_i_31,
	freq_mod_i_16,
	phi_inc_i_16,
	freq_mod_i_17,
	phi_inc_i_17,
	freq_mod_i_18,
	phi_inc_i_18,
	freq_mod_i_19,
	phi_inc_i_19,
	freq_mod_i_20,
	phi_inc_i_20,
	freq_mod_i_21,
	phi_inc_i_21,
	freq_mod_i_22,
	phi_inc_i_22,
	freq_mod_i_23,
	phi_inc_i_23,
	freq_mod_i_15,
	phi_inc_i_15,
	freq_mod_i_14,
	phi_inc_i_14,
	freq_mod_i_13,
	phi_inc_i_13,
	freq_mod_i_12,
	phi_inc_i_12,
	freq_mod_i_11,
	phi_inc_i_11,
	freq_mod_i_10,
	phi_inc_i_10,
	freq_mod_i_9,
	phi_inc_i_9,
	freq_mod_i_8,
	phi_inc_i_8,
	freq_mod_i_7,
	phi_inc_i_7,
	freq_mod_i_6,
	phi_inc_i_6,
	freq_mod_i_5,
	phi_inc_i_5,
	freq_mod_i_4,
	phi_inc_i_4,
	freq_mod_i_3,
	phi_inc_i_3,
	freq_mod_i_2,
	phi_inc_i_2,
	freq_mod_i_1,
	phi_inc_i_1,
	freq_mod_i_0,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	data_ready;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
input 	GND_port;
input 	NJQG9082;
input 	clk;
input 	clken;
input 	reset_n;
input 	phase_mod_i_8;
input 	phase_mod_i_9;
input 	phase_mod_i_10;
input 	phase_mod_i_11;
input 	phase_mod_i_12;
input 	phase_mod_i_13;
input 	phase_mod_i_14;
input 	phase_mod_i_15;
input 	phase_mod_i_0;
input 	phase_mod_i_1;
input 	phase_mod_i_2;
input 	phase_mod_i_3;
input 	phase_mod_i_4;
input 	phase_mod_i_5;
input 	phase_mod_i_6;
input 	phase_mod_i_7;
input 	freq_mod_i_24;
input 	phi_inc_i_24;
input 	freq_mod_i_25;
input 	phi_inc_i_25;
input 	freq_mod_i_26;
input 	phi_inc_i_26;
input 	freq_mod_i_27;
input 	phi_inc_i_27;
input 	freq_mod_i_28;
input 	phi_inc_i_28;
input 	freq_mod_i_29;
input 	phi_inc_i_29;
input 	freq_mod_i_30;
input 	phi_inc_i_30;
input 	freq_mod_i_31;
input 	phi_inc_i_31;
input 	freq_mod_i_16;
input 	phi_inc_i_16;
input 	freq_mod_i_17;
input 	phi_inc_i_17;
input 	freq_mod_i_18;
input 	phi_inc_i_18;
input 	freq_mod_i_19;
input 	phi_inc_i_19;
input 	freq_mod_i_20;
input 	phi_inc_i_20;
input 	freq_mod_i_21;
input 	phi_inc_i_21;
input 	freq_mod_i_22;
input 	phi_inc_i_22;
input 	freq_mod_i_23;
input 	phi_inc_i_23;
input 	freq_mod_i_15;
input 	phi_inc_i_15;
input 	freq_mod_i_14;
input 	phi_inc_i_14;
input 	freq_mod_i_13;
input 	phi_inc_i_13;
input 	freq_mod_i_12;
input 	phi_inc_i_12;
input 	freq_mod_i_11;
input 	phi_inc_i_11;
input 	freq_mod_i_10;
input 	phi_inc_i_10;
input 	freq_mod_i_9;
input 	phi_inc_i_9;
input 	freq_mod_i_8;
input 	phi_inc_i_8;
input 	freq_mod_i_7;
input 	phi_inc_i_7;
input 	freq_mod_i_6;
input 	phi_inc_i_6;
input 	freq_mod_i_5;
input 	phi_inc_i_5;
input 	freq_mod_i_4;
input 	phi_inc_i_4;
input 	freq_mod_i_3;
input 	phi_inc_i_3;
input 	freq_mod_i_2;
input 	phi_inc_i_2;
input 	freq_mod_i_1;
input 	phi_inc_i_1;
input 	freq_mod_i_0;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ux0220|altsyncram_component|auto_generated|q_a[0] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[0] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[1] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[1] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[2] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[2] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[3] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[3] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[4] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[4] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[5] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[5] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[6] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[6] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[7] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[7] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[8] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[8] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[9] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[9] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[10] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[10] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[11] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[11] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[12] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[12] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[13] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[13] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[14] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[14] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[15] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[15] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[16] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[16] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[17] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[17] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[18] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[18] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[19] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[19] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[20] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[20] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[21] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[21] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[22] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[22] ;
wire \ux0220|altsyncram_component|auto_generated|q_a[23] ;
wire \ux0220|altsyncram_component|auto_generated|q_b[23] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[0] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[1] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[2] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[3] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[4] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[5] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[6] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[7] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[8] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[9] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[10] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[11] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[12] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[13] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[14] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[15] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[16] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[17] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[18] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[19] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[20] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[21] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[22] ;
wire \ux0123|altsyncram_component0|auto_generated|q_a[23] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[0] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[1] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[2] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[3] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[4] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[5] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[6] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[7] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[8] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[9] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[10] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[11] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[12] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[13] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[14] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[15] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[16] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[17] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[18] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[19] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[20] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[21] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[22] ;
wire \ux0122|altsyncram_component0|auto_generated|q_a[23] ;
wire \ux008|rom_add_cc_temp[0]~q ;
wire \ux008|rom_add_cc_temp[1]~q ;
wire \ux008|rom_add_cc_temp[2]~q ;
wire \ux008|rom_add_cc_temp[3]~q ;
wire \ux008|rom_add_cc_temp[4]~q ;
wire \ux008|rom_add_cc_temp[5]~q ;
wire \ux008|rom_add_cs[6]~q ;
wire \ux008|rom_add_cs[7]~q ;
wire \ux008|rom_add_cc_temp[6]~q ;
wire \ux008|rom_add_cc_temp[7]~q ;
wire \ux008|rom_add_f[0]~q ;
wire \ux008|rom_add_f[1]~q ;
wire \ux008|rom_add_f[2]~q ;
wire \ux008|rom_add_f[3]~q ;
wire \ux008|rom_add_f[4]~q ;
wire \ux008|rom_add_f[5]~q ;
wire \ux008|rom_add_f[6]~q ;
wire \ux008|rom_add_f[7]~q ;
wire \ux002|dxxpdo[13]~q ;
wire \ux002|dxxpdo[14]~q ;
wire \ux002|dxxpdo[15]~q ;
wire \ux002|dxxpdo[16]~q ;
wire \ux002|dxxpdo[17]~q ;
wire \ux002|dxxpdo[18]~q ;
wire \ux002|dxxpdo[19]~q ;
wire \ux002|dxxpdo[20]~q ;
wire \ux002|dxxpdo[5]~q ;
wire \ux002|dxxpdo[6]~q ;
wire \ux002|dxxpdo[7]~q ;
wire \ux002|dxxpdo[8]~q ;
wire \ux002|dxxpdo[9]~q ;
wire \ux002|dxxpdo[10]~q ;
wire \ux002|dxxpdo[11]~q ;
wire \ux002|dxxpdo[12]~q ;
wire \ux001|dxxrv[3]~q ;
wire \ux001|dxxrv[2]~q ;
wire \ux001|dxxrv[1]~q ;
wire \ux001|dxxrv[0]~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe47~q ;
wire \m0|result_a[28]~0_combout ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe24~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe35~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe48~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe25~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe26~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe27~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe28~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe29~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe30~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe31~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe32~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe33~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe34~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe36~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe37~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe38~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe39~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe40~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe41~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe42~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe43~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe44~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe45~q ;
wire \m0|a_0|lpm_add_sub_component|auto_generated|dffe46~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[8]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[9]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[10]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[11]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[12]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[13]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[14]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[15]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[0]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[1]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[2]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[3]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[4]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[5]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[6]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[7]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[24]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[25]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[26]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[27]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[28]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[29]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[30]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[31]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[16]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[17]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[18]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[19]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[20]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[21]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[22]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[23]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[15]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[14]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[24]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[25]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[26]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[27]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[28]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[29]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[30]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[31]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[16]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[13]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[17]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[18]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[19]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[20]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[21]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[22]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[23]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[15]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[12]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[14]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[11]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[13]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[12]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[11]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[10]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[9]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[8]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[7]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[6]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[5]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[4]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[3]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[2]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[1]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[0]~q ;


sine_asj_dxx ux002(
	.dxxpdo_13(\ux002|dxxpdo[13]~q ),
	.dxxpdo_14(\ux002|dxxpdo[14]~q ),
	.dxxpdo_15(\ux002|dxxpdo[15]~q ),
	.dxxpdo_16(\ux002|dxxpdo[16]~q ),
	.dxxpdo_17(\ux002|dxxpdo[17]~q ),
	.dxxpdo_18(\ux002|dxxpdo[18]~q ),
	.dxxpdo_19(\ux002|dxxpdo[19]~q ),
	.dxxpdo_20(\ux002|dxxpdo[20]~q ),
	.dxxpdo_5(\ux002|dxxpdo[5]~q ),
	.dxxpdo_6(\ux002|dxxpdo[6]~q ),
	.dxxpdo_7(\ux002|dxxpdo[7]~q ),
	.dxxpdo_8(\ux002|dxxpdo[8]~q ),
	.dxxpdo_9(\ux002|dxxpdo[9]~q ),
	.dxxpdo_10(\ux002|dxxpdo[10]~q ),
	.dxxpdo_11(\ux002|dxxpdo[11]~q ),
	.dxxpdo_12(\ux002|dxxpdo[12]~q ),
	.dxxrv_3(\ux001|dxxrv[3]~q ),
	.dxxrv_2(\ux001|dxxrv[2]~q ),
	.dxxrv_1(\ux001|dxxrv[1]~q ),
	.dxxrv_0(\ux001|dxxrv[0]~q ),
	.result_a_28(\m0|result_a[28]~0_combout ),
	.pipeline_dffe_24(\ux000|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_25(\ux000|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_26(\ux000|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_27(\ux000|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_28(\ux000|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_29(\ux000|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_30(\ux000|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_31(\ux000|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_16(\ux000|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\ux000|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\ux000|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_19(\ux000|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_20(\ux000|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_21(\ux000|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_22(\ux000|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_23(\ux000|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_15(\ux000|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_14(\ux000|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\ux000|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_12(\ux000|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\ux000|acc|auto_generated|pipeline_dffe[11]~q ),
	.NJQG9082(NJQG9082),
	.clk(clk),
	.reset_n(reset_n));

sine_asj_dxx_g ux001(
	.dxxrv_3(\ux001|dxxrv[3]~q ),
	.dxxrv_2(\ux001|dxxrv[2]~q ),
	.dxxrv_1(\ux001|dxxrv[1]~q ),
	.dxxrv_0(\ux001|dxxrv[0]~q ),
	.result_a_28(\m0|result_a[28]~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

sine_asj_altqmcpipe ux000(
	.result_a_28(\m0|result_a[28]~0_combout ),
	.pipeline_dffe_24(\ux000|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_25(\ux000|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_26(\ux000|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_27(\ux000|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_28(\ux000|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_29(\ux000|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_30(\ux000|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_31(\ux000|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_16(\ux000|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\ux000|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\ux000|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_19(\ux000|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_20(\ux000|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_21(\ux000|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_22(\ux000|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_23(\ux000|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_15(\ux000|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_14(\ux000|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_241(\ux003|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_251(\ux003|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_261(\ux003|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_271(\ux003|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_281(\ux003|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_291(\ux003|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_301(\ux003|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_311(\ux003|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_161(\ux003|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_13(\ux000|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_171(\ux003|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_181(\ux003|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_191(\ux003|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_201(\ux003|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_211(\ux003|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_221(\ux003|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_231(\ux003|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_151(\ux003|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\ux000|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_141(\ux003|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_11(\ux000|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_131(\ux003|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_121(\ux003|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_111(\ux003|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\ux003|acc|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_9(\ux003|acc|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\ux003|acc|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\ux003|acc|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_6(\ux003|acc|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\ux003|acc|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\ux003|acc|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\ux003|acc|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\ux003|acc|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_1(\ux003|acc|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_0(\ux003|acc|auto_generated|pipeline_dffe[0]~q ),
	.clk(clk),
	.clken(clken),
	.reset_n(reset_n));

sine_asj_nco_mob_w blk0(
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.dffe47(\m0|a_0|lpm_add_sub_component|auto_generated|dffe47~q ),
	.result_a_28(\m0|result_a[28]~0_combout ),
	.dffe24(\m0|a_0|lpm_add_sub_component|auto_generated|dffe24~q ),
	.dffe35(\m0|a_0|lpm_add_sub_component|auto_generated|dffe35~q ),
	.dffe48(\m0|a_0|lpm_add_sub_component|auto_generated|dffe48~q ),
	.dffe25(\m0|a_0|lpm_add_sub_component|auto_generated|dffe25~q ),
	.dffe26(\m0|a_0|lpm_add_sub_component|auto_generated|dffe26~q ),
	.dffe27(\m0|a_0|lpm_add_sub_component|auto_generated|dffe27~q ),
	.dffe28(\m0|a_0|lpm_add_sub_component|auto_generated|dffe28~q ),
	.dffe29(\m0|a_0|lpm_add_sub_component|auto_generated|dffe29~q ),
	.dffe30(\m0|a_0|lpm_add_sub_component|auto_generated|dffe30~q ),
	.dffe31(\m0|a_0|lpm_add_sub_component|auto_generated|dffe31~q ),
	.dffe32(\m0|a_0|lpm_add_sub_component|auto_generated|dffe32~q ),
	.dffe33(\m0|a_0|lpm_add_sub_component|auto_generated|dffe33~q ),
	.dffe34(\m0|a_0|lpm_add_sub_component|auto_generated|dffe34~q ),
	.dffe36(\m0|a_0|lpm_add_sub_component|auto_generated|dffe36~q ),
	.dffe37(\m0|a_0|lpm_add_sub_component|auto_generated|dffe37~q ),
	.dffe38(\m0|a_0|lpm_add_sub_component|auto_generated|dffe38~q ),
	.dffe39(\m0|a_0|lpm_add_sub_component|auto_generated|dffe39~q ),
	.dffe40(\m0|a_0|lpm_add_sub_component|auto_generated|dffe40~q ),
	.dffe41(\m0|a_0|lpm_add_sub_component|auto_generated|dffe41~q ),
	.dffe42(\m0|a_0|lpm_add_sub_component|auto_generated|dffe42~q ),
	.dffe43(\m0|a_0|lpm_add_sub_component|auto_generated|dffe43~q ),
	.dffe44(\m0|a_0|lpm_add_sub_component|auto_generated|dffe44~q ),
	.dffe45(\m0|a_0|lpm_add_sub_component|auto_generated|dffe45~q ),
	.dffe46(\m0|a_0|lpm_add_sub_component|auto_generated|dffe46~q ),
	.clk(clk),
	.clken(clken),
	.reset_n(reset_n));

sine_mac_i_lpmd m0(
	.q_a_0(\ux0220|altsyncram_component|auto_generated|q_a[0] ),
	.q_b_0(\ux0220|altsyncram_component|auto_generated|q_b[0] ),
	.q_a_1(\ux0220|altsyncram_component|auto_generated|q_a[1] ),
	.q_b_1(\ux0220|altsyncram_component|auto_generated|q_b[1] ),
	.q_a_2(\ux0220|altsyncram_component|auto_generated|q_a[2] ),
	.q_b_2(\ux0220|altsyncram_component|auto_generated|q_b[2] ),
	.q_a_3(\ux0220|altsyncram_component|auto_generated|q_a[3] ),
	.q_b_3(\ux0220|altsyncram_component|auto_generated|q_b[3] ),
	.q_a_4(\ux0220|altsyncram_component|auto_generated|q_a[4] ),
	.q_b_4(\ux0220|altsyncram_component|auto_generated|q_b[4] ),
	.q_a_5(\ux0220|altsyncram_component|auto_generated|q_a[5] ),
	.q_b_5(\ux0220|altsyncram_component|auto_generated|q_b[5] ),
	.q_a_6(\ux0220|altsyncram_component|auto_generated|q_a[6] ),
	.q_b_6(\ux0220|altsyncram_component|auto_generated|q_b[6] ),
	.q_a_7(\ux0220|altsyncram_component|auto_generated|q_a[7] ),
	.q_b_7(\ux0220|altsyncram_component|auto_generated|q_b[7] ),
	.q_a_8(\ux0220|altsyncram_component|auto_generated|q_a[8] ),
	.q_b_8(\ux0220|altsyncram_component|auto_generated|q_b[8] ),
	.q_a_9(\ux0220|altsyncram_component|auto_generated|q_a[9] ),
	.q_b_9(\ux0220|altsyncram_component|auto_generated|q_b[9] ),
	.q_a_10(\ux0220|altsyncram_component|auto_generated|q_a[10] ),
	.q_b_10(\ux0220|altsyncram_component|auto_generated|q_b[10] ),
	.q_a_11(\ux0220|altsyncram_component|auto_generated|q_a[11] ),
	.q_b_11(\ux0220|altsyncram_component|auto_generated|q_b[11] ),
	.q_a_12(\ux0220|altsyncram_component|auto_generated|q_a[12] ),
	.q_b_12(\ux0220|altsyncram_component|auto_generated|q_b[12] ),
	.q_a_13(\ux0220|altsyncram_component|auto_generated|q_a[13] ),
	.q_b_13(\ux0220|altsyncram_component|auto_generated|q_b[13] ),
	.q_a_14(\ux0220|altsyncram_component|auto_generated|q_a[14] ),
	.q_b_14(\ux0220|altsyncram_component|auto_generated|q_b[14] ),
	.q_a_15(\ux0220|altsyncram_component|auto_generated|q_a[15] ),
	.q_b_15(\ux0220|altsyncram_component|auto_generated|q_b[15] ),
	.q_a_16(\ux0220|altsyncram_component|auto_generated|q_a[16] ),
	.q_b_16(\ux0220|altsyncram_component|auto_generated|q_b[16] ),
	.q_a_17(\ux0220|altsyncram_component|auto_generated|q_a[17] ),
	.q_b_17(\ux0220|altsyncram_component|auto_generated|q_b[17] ),
	.q_a_18(\ux0220|altsyncram_component|auto_generated|q_a[18] ),
	.q_b_18(\ux0220|altsyncram_component|auto_generated|q_b[18] ),
	.q_a_19(\ux0220|altsyncram_component|auto_generated|q_a[19] ),
	.q_b_19(\ux0220|altsyncram_component|auto_generated|q_b[19] ),
	.q_a_20(\ux0220|altsyncram_component|auto_generated|q_a[20] ),
	.q_b_20(\ux0220|altsyncram_component|auto_generated|q_b[20] ),
	.q_a_21(\ux0220|altsyncram_component|auto_generated|q_a[21] ),
	.q_b_21(\ux0220|altsyncram_component|auto_generated|q_b[21] ),
	.q_a_22(\ux0220|altsyncram_component|auto_generated|q_a[22] ),
	.q_b_22(\ux0220|altsyncram_component|auto_generated|q_b[22] ),
	.q_a_23(\ux0220|altsyncram_component|auto_generated|q_a[23] ),
	.q_b_23(\ux0220|altsyncram_component|auto_generated|q_b[23] ),
	.q_a_01(\ux0123|altsyncram_component0|auto_generated|q_a[0] ),
	.q_a_110(\ux0123|altsyncram_component0|auto_generated|q_a[1] ),
	.q_a_24(\ux0123|altsyncram_component0|auto_generated|q_a[2] ),
	.q_a_31(\ux0123|altsyncram_component0|auto_generated|q_a[3] ),
	.q_a_41(\ux0123|altsyncram_component0|auto_generated|q_a[4] ),
	.q_a_51(\ux0123|altsyncram_component0|auto_generated|q_a[5] ),
	.q_a_61(\ux0123|altsyncram_component0|auto_generated|q_a[6] ),
	.q_a_71(\ux0123|altsyncram_component0|auto_generated|q_a[7] ),
	.q_a_81(\ux0123|altsyncram_component0|auto_generated|q_a[8] ),
	.q_a_91(\ux0123|altsyncram_component0|auto_generated|q_a[9] ),
	.q_a_101(\ux0123|altsyncram_component0|auto_generated|q_a[10] ),
	.q_a_111(\ux0123|altsyncram_component0|auto_generated|q_a[11] ),
	.q_a_121(\ux0123|altsyncram_component0|auto_generated|q_a[12] ),
	.q_a_131(\ux0123|altsyncram_component0|auto_generated|q_a[13] ),
	.q_a_141(\ux0123|altsyncram_component0|auto_generated|q_a[14] ),
	.q_a_151(\ux0123|altsyncram_component0|auto_generated|q_a[15] ),
	.q_a_161(\ux0123|altsyncram_component0|auto_generated|q_a[16] ),
	.q_a_171(\ux0123|altsyncram_component0|auto_generated|q_a[17] ),
	.q_a_181(\ux0123|altsyncram_component0|auto_generated|q_a[18] ),
	.q_a_191(\ux0123|altsyncram_component0|auto_generated|q_a[19] ),
	.q_a_201(\ux0123|altsyncram_component0|auto_generated|q_a[20] ),
	.q_a_211(\ux0123|altsyncram_component0|auto_generated|q_a[21] ),
	.q_a_221(\ux0123|altsyncram_component0|auto_generated|q_a[22] ),
	.q_a_231(\ux0123|altsyncram_component0|auto_generated|q_a[23] ),
	.q_a_02(\ux0122|altsyncram_component0|auto_generated|q_a[0] ),
	.q_a_112(\ux0122|altsyncram_component0|auto_generated|q_a[1] ),
	.q_a_25(\ux0122|altsyncram_component0|auto_generated|q_a[2] ),
	.q_a_32(\ux0122|altsyncram_component0|auto_generated|q_a[3] ),
	.q_a_42(\ux0122|altsyncram_component0|auto_generated|q_a[4] ),
	.q_a_52(\ux0122|altsyncram_component0|auto_generated|q_a[5] ),
	.q_a_62(\ux0122|altsyncram_component0|auto_generated|q_a[6] ),
	.q_a_72(\ux0122|altsyncram_component0|auto_generated|q_a[7] ),
	.q_a_82(\ux0122|altsyncram_component0|auto_generated|q_a[8] ),
	.q_a_92(\ux0122|altsyncram_component0|auto_generated|q_a[9] ),
	.q_a_102(\ux0122|altsyncram_component0|auto_generated|q_a[10] ),
	.q_a_113(\ux0122|altsyncram_component0|auto_generated|q_a[11] ),
	.q_a_122(\ux0122|altsyncram_component0|auto_generated|q_a[12] ),
	.q_a_132(\ux0122|altsyncram_component0|auto_generated|q_a[13] ),
	.q_a_142(\ux0122|altsyncram_component0|auto_generated|q_a[14] ),
	.q_a_152(\ux0122|altsyncram_component0|auto_generated|q_a[15] ),
	.q_a_162(\ux0122|altsyncram_component0|auto_generated|q_a[16] ),
	.q_a_172(\ux0122|altsyncram_component0|auto_generated|q_a[17] ),
	.q_a_182(\ux0122|altsyncram_component0|auto_generated|q_a[18] ),
	.q_a_192(\ux0122|altsyncram_component0|auto_generated|q_a[19] ),
	.q_a_202(\ux0122|altsyncram_component0|auto_generated|q_a[20] ),
	.q_a_212(\ux0122|altsyncram_component0|auto_generated|q_a[21] ),
	.q_a_222(\ux0122|altsyncram_component0|auto_generated|q_a[22] ),
	.q_a_232(\ux0122|altsyncram_component0|auto_generated|q_a[23] ),
	.dffe47(\m0|a_0|lpm_add_sub_component|auto_generated|dffe47~q ),
	.result_a_28(\m0|result_a[28]~0_combout ),
	.dffe24(\m0|a_0|lpm_add_sub_component|auto_generated|dffe24~q ),
	.dffe35(\m0|a_0|lpm_add_sub_component|auto_generated|dffe35~q ),
	.dffe48(\m0|a_0|lpm_add_sub_component|auto_generated|dffe48~q ),
	.dffe25(\m0|a_0|lpm_add_sub_component|auto_generated|dffe25~q ),
	.dffe26(\m0|a_0|lpm_add_sub_component|auto_generated|dffe26~q ),
	.dffe27(\m0|a_0|lpm_add_sub_component|auto_generated|dffe27~q ),
	.dffe28(\m0|a_0|lpm_add_sub_component|auto_generated|dffe28~q ),
	.dffe29(\m0|a_0|lpm_add_sub_component|auto_generated|dffe29~q ),
	.dffe30(\m0|a_0|lpm_add_sub_component|auto_generated|dffe30~q ),
	.dffe31(\m0|a_0|lpm_add_sub_component|auto_generated|dffe31~q ),
	.dffe32(\m0|a_0|lpm_add_sub_component|auto_generated|dffe32~q ),
	.dffe33(\m0|a_0|lpm_add_sub_component|auto_generated|dffe33~q ),
	.dffe34(\m0|a_0|lpm_add_sub_component|auto_generated|dffe34~q ),
	.dffe36(\m0|a_0|lpm_add_sub_component|auto_generated|dffe36~q ),
	.dffe37(\m0|a_0|lpm_add_sub_component|auto_generated|dffe37~q ),
	.dffe38(\m0|a_0|lpm_add_sub_component|auto_generated|dffe38~q ),
	.dffe39(\m0|a_0|lpm_add_sub_component|auto_generated|dffe39~q ),
	.dffe40(\m0|a_0|lpm_add_sub_component|auto_generated|dffe40~q ),
	.dffe41(\m0|a_0|lpm_add_sub_component|auto_generated|dffe41~q ),
	.dffe42(\m0|a_0|lpm_add_sub_component|auto_generated|dffe42~q ),
	.dffe43(\m0|a_0|lpm_add_sub_component|auto_generated|dffe43~q ),
	.dffe44(\m0|a_0|lpm_add_sub_component|auto_generated|dffe44~q ),
	.dffe45(\m0|a_0|lpm_add_sub_component|auto_generated|dffe45~q ),
	.dffe46(\m0|a_0|lpm_add_sub_component|auto_generated|dffe46~q ),
	.clk(clk),
	.clken(clken),
	.reset_n(reset_n));

sine_asj_nco_as_m_cen_1 ux0123(
	.q_a_0(\ux0123|altsyncram_component0|auto_generated|q_a[0] ),
	.q_a_1(\ux0123|altsyncram_component0|auto_generated|q_a[1] ),
	.q_a_2(\ux0123|altsyncram_component0|auto_generated|q_a[2] ),
	.q_a_3(\ux0123|altsyncram_component0|auto_generated|q_a[3] ),
	.q_a_4(\ux0123|altsyncram_component0|auto_generated|q_a[4] ),
	.q_a_5(\ux0123|altsyncram_component0|auto_generated|q_a[5] ),
	.q_a_6(\ux0123|altsyncram_component0|auto_generated|q_a[6] ),
	.q_a_7(\ux0123|altsyncram_component0|auto_generated|q_a[7] ),
	.q_a_8(\ux0123|altsyncram_component0|auto_generated|q_a[8] ),
	.q_a_9(\ux0123|altsyncram_component0|auto_generated|q_a[9] ),
	.q_a_10(\ux0123|altsyncram_component0|auto_generated|q_a[10] ),
	.q_a_11(\ux0123|altsyncram_component0|auto_generated|q_a[11] ),
	.q_a_12(\ux0123|altsyncram_component0|auto_generated|q_a[12] ),
	.q_a_13(\ux0123|altsyncram_component0|auto_generated|q_a[13] ),
	.q_a_14(\ux0123|altsyncram_component0|auto_generated|q_a[14] ),
	.q_a_15(\ux0123|altsyncram_component0|auto_generated|q_a[15] ),
	.q_a_16(\ux0123|altsyncram_component0|auto_generated|q_a[16] ),
	.q_a_17(\ux0123|altsyncram_component0|auto_generated|q_a[17] ),
	.q_a_18(\ux0123|altsyncram_component0|auto_generated|q_a[18] ),
	.q_a_19(\ux0123|altsyncram_component0|auto_generated|q_a[19] ),
	.q_a_20(\ux0123|altsyncram_component0|auto_generated|q_a[20] ),
	.q_a_21(\ux0123|altsyncram_component0|auto_generated|q_a[21] ),
	.q_a_22(\ux0123|altsyncram_component0|auto_generated|q_a[22] ),
	.q_a_23(\ux0123|altsyncram_component0|auto_generated|q_a[23] ),
	.rom_add_f_0(\ux008|rom_add_f[0]~q ),
	.rom_add_f_1(\ux008|rom_add_f[1]~q ),
	.rom_add_f_2(\ux008|rom_add_f[2]~q ),
	.rom_add_f_3(\ux008|rom_add_f[3]~q ),
	.rom_add_f_4(\ux008|rom_add_f[4]~q ),
	.rom_add_f_5(\ux008|rom_add_f[5]~q ),
	.rom_add_f_6(\ux008|rom_add_f[6]~q ),
	.rom_add_f_7(\ux008|rom_add_f[7]~q ),
	.clk(clk),
	.clken(clken));

sine_asj_nco_as_m_cen ux0122(
	.q_a_0(\ux0122|altsyncram_component0|auto_generated|q_a[0] ),
	.q_a_1(\ux0122|altsyncram_component0|auto_generated|q_a[1] ),
	.q_a_2(\ux0122|altsyncram_component0|auto_generated|q_a[2] ),
	.q_a_3(\ux0122|altsyncram_component0|auto_generated|q_a[3] ),
	.q_a_4(\ux0122|altsyncram_component0|auto_generated|q_a[4] ),
	.q_a_5(\ux0122|altsyncram_component0|auto_generated|q_a[5] ),
	.q_a_6(\ux0122|altsyncram_component0|auto_generated|q_a[6] ),
	.q_a_7(\ux0122|altsyncram_component0|auto_generated|q_a[7] ),
	.q_a_8(\ux0122|altsyncram_component0|auto_generated|q_a[8] ),
	.q_a_9(\ux0122|altsyncram_component0|auto_generated|q_a[9] ),
	.q_a_10(\ux0122|altsyncram_component0|auto_generated|q_a[10] ),
	.q_a_11(\ux0122|altsyncram_component0|auto_generated|q_a[11] ),
	.q_a_12(\ux0122|altsyncram_component0|auto_generated|q_a[12] ),
	.q_a_13(\ux0122|altsyncram_component0|auto_generated|q_a[13] ),
	.q_a_14(\ux0122|altsyncram_component0|auto_generated|q_a[14] ),
	.q_a_15(\ux0122|altsyncram_component0|auto_generated|q_a[15] ),
	.q_a_16(\ux0122|altsyncram_component0|auto_generated|q_a[16] ),
	.q_a_17(\ux0122|altsyncram_component0|auto_generated|q_a[17] ),
	.q_a_18(\ux0122|altsyncram_component0|auto_generated|q_a[18] ),
	.q_a_19(\ux0122|altsyncram_component0|auto_generated|q_a[19] ),
	.q_a_20(\ux0122|altsyncram_component0|auto_generated|q_a[20] ),
	.q_a_21(\ux0122|altsyncram_component0|auto_generated|q_a[21] ),
	.q_a_22(\ux0122|altsyncram_component0|auto_generated|q_a[22] ),
	.q_a_23(\ux0122|altsyncram_component0|auto_generated|q_a[23] ),
	.rom_add_f_0(\ux008|rom_add_f[0]~q ),
	.rom_add_f_1(\ux008|rom_add_f[1]~q ),
	.rom_add_f_2(\ux008|rom_add_f[2]~q ),
	.rom_add_f_3(\ux008|rom_add_f[3]~q ),
	.rom_add_f_4(\ux008|rom_add_f[4]~q ),
	.rom_add_f_5(\ux008|rom_add_f[5]~q ),
	.rom_add_f_6(\ux008|rom_add_f[6]~q ),
	.rom_add_f_7(\ux008|rom_add_f[7]~q ),
	.clk(clk),
	.clken(clken));

sine_asj_nco_as_m_dp_cen ux0220(
	.q_a_0(\ux0220|altsyncram_component|auto_generated|q_a[0] ),
	.q_b_0(\ux0220|altsyncram_component|auto_generated|q_b[0] ),
	.q_a_1(\ux0220|altsyncram_component|auto_generated|q_a[1] ),
	.q_b_1(\ux0220|altsyncram_component|auto_generated|q_b[1] ),
	.q_a_2(\ux0220|altsyncram_component|auto_generated|q_a[2] ),
	.q_b_2(\ux0220|altsyncram_component|auto_generated|q_b[2] ),
	.q_a_3(\ux0220|altsyncram_component|auto_generated|q_a[3] ),
	.q_b_3(\ux0220|altsyncram_component|auto_generated|q_b[3] ),
	.q_a_4(\ux0220|altsyncram_component|auto_generated|q_a[4] ),
	.q_b_4(\ux0220|altsyncram_component|auto_generated|q_b[4] ),
	.q_a_5(\ux0220|altsyncram_component|auto_generated|q_a[5] ),
	.q_b_5(\ux0220|altsyncram_component|auto_generated|q_b[5] ),
	.q_a_6(\ux0220|altsyncram_component|auto_generated|q_a[6] ),
	.q_b_6(\ux0220|altsyncram_component|auto_generated|q_b[6] ),
	.q_a_7(\ux0220|altsyncram_component|auto_generated|q_a[7] ),
	.q_b_7(\ux0220|altsyncram_component|auto_generated|q_b[7] ),
	.q_a_8(\ux0220|altsyncram_component|auto_generated|q_a[8] ),
	.q_b_8(\ux0220|altsyncram_component|auto_generated|q_b[8] ),
	.q_a_9(\ux0220|altsyncram_component|auto_generated|q_a[9] ),
	.q_b_9(\ux0220|altsyncram_component|auto_generated|q_b[9] ),
	.q_a_10(\ux0220|altsyncram_component|auto_generated|q_a[10] ),
	.q_b_10(\ux0220|altsyncram_component|auto_generated|q_b[10] ),
	.q_a_11(\ux0220|altsyncram_component|auto_generated|q_a[11] ),
	.q_b_11(\ux0220|altsyncram_component|auto_generated|q_b[11] ),
	.q_a_12(\ux0220|altsyncram_component|auto_generated|q_a[12] ),
	.q_b_12(\ux0220|altsyncram_component|auto_generated|q_b[12] ),
	.q_a_13(\ux0220|altsyncram_component|auto_generated|q_a[13] ),
	.q_b_13(\ux0220|altsyncram_component|auto_generated|q_b[13] ),
	.q_a_14(\ux0220|altsyncram_component|auto_generated|q_a[14] ),
	.q_b_14(\ux0220|altsyncram_component|auto_generated|q_b[14] ),
	.q_a_15(\ux0220|altsyncram_component|auto_generated|q_a[15] ),
	.q_b_15(\ux0220|altsyncram_component|auto_generated|q_b[15] ),
	.q_a_16(\ux0220|altsyncram_component|auto_generated|q_a[16] ),
	.q_b_16(\ux0220|altsyncram_component|auto_generated|q_b[16] ),
	.q_a_17(\ux0220|altsyncram_component|auto_generated|q_a[17] ),
	.q_b_17(\ux0220|altsyncram_component|auto_generated|q_b[17] ),
	.q_a_18(\ux0220|altsyncram_component|auto_generated|q_a[18] ),
	.q_b_18(\ux0220|altsyncram_component|auto_generated|q_b[18] ),
	.q_a_19(\ux0220|altsyncram_component|auto_generated|q_a[19] ),
	.q_b_19(\ux0220|altsyncram_component|auto_generated|q_b[19] ),
	.q_a_20(\ux0220|altsyncram_component|auto_generated|q_a[20] ),
	.q_b_20(\ux0220|altsyncram_component|auto_generated|q_b[20] ),
	.q_a_21(\ux0220|altsyncram_component|auto_generated|q_a[21] ),
	.q_b_21(\ux0220|altsyncram_component|auto_generated|q_b[21] ),
	.q_a_22(\ux0220|altsyncram_component|auto_generated|q_a[22] ),
	.q_b_22(\ux0220|altsyncram_component|auto_generated|q_b[22] ),
	.q_a_23(\ux0220|altsyncram_component|auto_generated|q_a[23] ),
	.q_b_23(\ux0220|altsyncram_component|auto_generated|q_b[23] ),
	.rom_add_cc_temp_0(\ux008|rom_add_cc_temp[0]~q ),
	.rom_add_cc_temp_1(\ux008|rom_add_cc_temp[1]~q ),
	.rom_add_cc_temp_2(\ux008|rom_add_cc_temp[2]~q ),
	.rom_add_cc_temp_3(\ux008|rom_add_cc_temp[3]~q ),
	.rom_add_cc_temp_4(\ux008|rom_add_cc_temp[4]~q ),
	.rom_add_cc_temp_5(\ux008|rom_add_cc_temp[5]~q ),
	.rom_add_cs_6(\ux008|rom_add_cs[6]~q ),
	.rom_add_cs_7(\ux008|rom_add_cs[7]~q ),
	.rom_add_cc_temp_6(\ux008|rom_add_cc_temp[6]~q ),
	.rom_add_cc_temp_7(\ux008|rom_add_cc_temp[7]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.clken(clken));

sine_asj_gam_dp ux008(
	.rom_add_cc_temp_0(\ux008|rom_add_cc_temp[0]~q ),
	.rom_add_cc_temp_1(\ux008|rom_add_cc_temp[1]~q ),
	.rom_add_cc_temp_2(\ux008|rom_add_cc_temp[2]~q ),
	.rom_add_cc_temp_3(\ux008|rom_add_cc_temp[3]~q ),
	.rom_add_cc_temp_4(\ux008|rom_add_cc_temp[4]~q ),
	.rom_add_cc_temp_5(\ux008|rom_add_cc_temp[5]~q ),
	.rom_add_cs_6(\ux008|rom_add_cs[6]~q ),
	.rom_add_cs_7(\ux008|rom_add_cs[7]~q ),
	.rom_add_cc_temp_6(\ux008|rom_add_cc_temp[6]~q ),
	.rom_add_cc_temp_7(\ux008|rom_add_cc_temp[7]~q ),
	.rom_add_f_0(\ux008|rom_add_f[0]~q ),
	.rom_add_f_1(\ux008|rom_add_f[1]~q ),
	.rom_add_f_2(\ux008|rom_add_f[2]~q ),
	.rom_add_f_3(\ux008|rom_add_f[3]~q ),
	.rom_add_f_4(\ux008|rom_add_f[4]~q ),
	.rom_add_f_5(\ux008|rom_add_f[5]~q ),
	.rom_add_f_6(\ux008|rom_add_f[6]~q ),
	.rom_add_f_7(\ux008|rom_add_f[7]~q ),
	.result_a_28(\m0|result_a[28]~0_combout ),
	.pipeline_dffe_8(\ux004|acc|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\ux004|acc|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\ux004|acc|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\ux004|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\ux004|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\ux004|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\ux004|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_15(\ux004|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_0(\ux004|acc|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\ux004|acc|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\ux004|acc|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\ux004|acc|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\ux004|acc|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\ux004|acc|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\ux004|acc|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\ux004|acc|auto_generated|pipeline_dffe[7]~q ),
	.clk(clk),
	.reset_n(reset_n));

sine_asj_nco_pxx ux004(
	.dxxpdo_13(\ux002|dxxpdo[13]~q ),
	.dxxpdo_14(\ux002|dxxpdo[14]~q ),
	.dxxpdo_15(\ux002|dxxpdo[15]~q ),
	.dxxpdo_16(\ux002|dxxpdo[16]~q ),
	.dxxpdo_17(\ux002|dxxpdo[17]~q ),
	.dxxpdo_18(\ux002|dxxpdo[18]~q ),
	.dxxpdo_19(\ux002|dxxpdo[19]~q ),
	.dxxpdo_20(\ux002|dxxpdo[20]~q ),
	.dxxpdo_5(\ux002|dxxpdo[5]~q ),
	.dxxpdo_6(\ux002|dxxpdo[6]~q ),
	.dxxpdo_7(\ux002|dxxpdo[7]~q ),
	.dxxpdo_8(\ux002|dxxpdo[8]~q ),
	.dxxpdo_9(\ux002|dxxpdo[9]~q ),
	.dxxpdo_10(\ux002|dxxpdo[10]~q ),
	.dxxpdo_11(\ux002|dxxpdo[11]~q ),
	.dxxpdo_12(\ux002|dxxpdo[12]~q ),
	.result_a_28(\m0|result_a[28]~0_combout ),
	.pipeline_dffe_8(\ux004|acc|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\ux004|acc|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\ux004|acc|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\ux004|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\ux004|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\ux004|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\ux004|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_15(\ux004|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_0(\ux004|acc|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\ux004|acc|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\ux004|acc|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\ux004|acc|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\ux004|acc|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\ux004|acc|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\ux004|acc|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\ux004|acc|auto_generated|pipeline_dffe[7]~q ),
	.clk(clk),
	.clken(clken),
	.reset_n(reset_n),
	.phase_mod_i_8(phase_mod_i_8),
	.phase_mod_i_9(phase_mod_i_9),
	.phase_mod_i_10(phase_mod_i_10),
	.phase_mod_i_11(phase_mod_i_11),
	.phase_mod_i_12(phase_mod_i_12),
	.phase_mod_i_13(phase_mod_i_13),
	.phase_mod_i_14(phase_mod_i_14),
	.phase_mod_i_15(phase_mod_i_15),
	.phase_mod_i_0(phase_mod_i_0),
	.phase_mod_i_1(phase_mod_i_1),
	.phase_mod_i_2(phase_mod_i_2),
	.phase_mod_i_3(phase_mod_i_3),
	.phase_mod_i_4(phase_mod_i_4),
	.phase_mod_i_5(phase_mod_i_5),
	.phase_mod_i_6(phase_mod_i_6),
	.phase_mod_i_7(phase_mod_i_7));

sine_asj_nco_fxx ux003(
	.pipeline_dffe_24(\ux003|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_25(\ux003|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_26(\ux003|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_27(\ux003|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_28(\ux003|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_29(\ux003|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_30(\ux003|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_31(\ux003|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_16(\ux003|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\ux003|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\ux003|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_19(\ux003|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_20(\ux003|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_21(\ux003|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_22(\ux003|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_23(\ux003|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_15(\ux003|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_14(\ux003|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\ux003|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_12(\ux003|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\ux003|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\ux003|acc|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_9(\ux003|acc|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\ux003|acc|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\ux003|acc|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_6(\ux003|acc|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\ux003|acc|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\ux003|acc|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\ux003|acc|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\ux003|acc|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_1(\ux003|acc|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_0(\ux003|acc|auto_generated|pipeline_dffe[0]~q ),
	.clk(clk),
	.clken(clken),
	.reset_n(reset_n),
	.freq_mod_i_24(freq_mod_i_24),
	.phi_inc_i_24(phi_inc_i_24),
	.freq_mod_i_25(freq_mod_i_25),
	.phi_inc_i_25(phi_inc_i_25),
	.freq_mod_i_26(freq_mod_i_26),
	.phi_inc_i_26(phi_inc_i_26),
	.freq_mod_i_27(freq_mod_i_27),
	.phi_inc_i_27(phi_inc_i_27),
	.freq_mod_i_28(freq_mod_i_28),
	.phi_inc_i_28(phi_inc_i_28),
	.freq_mod_i_29(freq_mod_i_29),
	.phi_inc_i_29(phi_inc_i_29),
	.freq_mod_i_30(freq_mod_i_30),
	.phi_inc_i_30(phi_inc_i_30),
	.freq_mod_i_31(freq_mod_i_31),
	.phi_inc_i_31(phi_inc_i_31),
	.freq_mod_i_16(freq_mod_i_16),
	.phi_inc_i_16(phi_inc_i_16),
	.freq_mod_i_17(freq_mod_i_17),
	.phi_inc_i_17(phi_inc_i_17),
	.freq_mod_i_18(freq_mod_i_18),
	.phi_inc_i_18(phi_inc_i_18),
	.freq_mod_i_19(freq_mod_i_19),
	.phi_inc_i_19(phi_inc_i_19),
	.freq_mod_i_20(freq_mod_i_20),
	.phi_inc_i_20(phi_inc_i_20),
	.freq_mod_i_21(freq_mod_i_21),
	.phi_inc_i_21(phi_inc_i_21),
	.freq_mod_i_22(freq_mod_i_22),
	.phi_inc_i_22(phi_inc_i_22),
	.freq_mod_i_23(freq_mod_i_23),
	.phi_inc_i_23(phi_inc_i_23),
	.freq_mod_i_15(freq_mod_i_15),
	.phi_inc_i_15(phi_inc_i_15),
	.freq_mod_i_14(freq_mod_i_14),
	.phi_inc_i_14(phi_inc_i_14),
	.freq_mod_i_13(freq_mod_i_13),
	.phi_inc_i_13(phi_inc_i_13),
	.freq_mod_i_12(freq_mod_i_12),
	.phi_inc_i_12(phi_inc_i_12),
	.freq_mod_i_11(freq_mod_i_11),
	.phi_inc_i_11(phi_inc_i_11),
	.freq_mod_i_10(freq_mod_i_10),
	.phi_inc_i_10(phi_inc_i_10),
	.freq_mod_i_9(freq_mod_i_9),
	.phi_inc_i_9(phi_inc_i_9),
	.freq_mod_i_8(freq_mod_i_8),
	.phi_inc_i_8(phi_inc_i_8),
	.freq_mod_i_7(freq_mod_i_7),
	.phi_inc_i_7(phi_inc_i_7),
	.freq_mod_i_6(freq_mod_i_6),
	.phi_inc_i_6(phi_inc_i_6),
	.freq_mod_i_5(freq_mod_i_5),
	.phi_inc_i_5(phi_inc_i_5),
	.freq_mod_i_4(freq_mod_i_4),
	.phi_inc_i_4(phi_inc_i_4),
	.freq_mod_i_3(freq_mod_i_3),
	.phi_inc_i_3(phi_inc_i_3),
	.freq_mod_i_2(freq_mod_i_2),
	.phi_inc_i_2(phi_inc_i_2),
	.freq_mod_i_1(freq_mod_i_1),
	.phi_inc_i_1(phi_inc_i_1),
	.freq_mod_i_0(freq_mod_i_0),
	.phi_inc_i_0(phi_inc_i_0));

sine_asj_nco_isdr ux710isdr(
	.data_ready1(data_ready),
	.clk(clk),
	.clken(clken),
	.reset_n(reset_n));

endmodule

module sine_asj_altqmcpipe (
	result_a_28,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_241,
	pipeline_dffe_251,
	pipeline_dffe_261,
	pipeline_dffe_271,
	pipeline_dffe_281,
	pipeline_dffe_291,
	pipeline_dffe_301,
	pipeline_dffe_311,
	pipeline_dffe_161,
	pipeline_dffe_13,
	pipeline_dffe_171,
	pipeline_dffe_181,
	pipeline_dffe_191,
	pipeline_dffe_201,
	pipeline_dffe_211,
	pipeline_dffe_221,
	pipeline_dffe_231,
	pipeline_dffe_151,
	pipeline_dffe_12,
	pipeline_dffe_141,
	pipeline_dffe_11,
	pipeline_dffe_131,
	pipeline_dffe_121,
	pipeline_dffe_111,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	clk,
	clken,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	result_a_28;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
input 	pipeline_dffe_241;
input 	pipeline_dffe_251;
input 	pipeline_dffe_261;
input 	pipeline_dffe_271;
input 	pipeline_dffe_281;
input 	pipeline_dffe_291;
input 	pipeline_dffe_301;
input 	pipeline_dffe_311;
input 	pipeline_dffe_161;
output 	pipeline_dffe_13;
input 	pipeline_dffe_171;
input 	pipeline_dffe_181;
input 	pipeline_dffe_191;
input 	pipeline_dffe_201;
input 	pipeline_dffe_211;
input 	pipeline_dffe_221;
input 	pipeline_dffe_231;
input 	pipeline_dffe_151;
output 	pipeline_dffe_12;
input 	pipeline_dffe_141;
output 	pipeline_dffe_11;
input 	pipeline_dffe_131;
input 	pipeline_dffe_121;
input 	pipeline_dffe_111;
input 	pipeline_dffe_10;
input 	pipeline_dffe_9;
input 	pipeline_dffe_8;
input 	pipeline_dffe_7;
input 	pipeline_dffe_6;
input 	pipeline_dffe_5;
input 	pipeline_dffe_4;
input 	pipeline_dffe_3;
input 	pipeline_dffe_2;
input 	pipeline_dffe_1;
input 	pipeline_dffe_0;
input 	clk;
input 	clken;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \phi_int_arr_reg[24]~q ;
wire \phi_int_arr_reg[25]~q ;
wire \phi_int_arr_reg[26]~q ;
wire \phi_int_arr_reg[27]~q ;
wire \phi_int_arr_reg[28]~q ;
wire \phi_int_arr_reg[29]~q ;
wire \phi_int_arr_reg[30]~q ;
wire \phi_int_arr_reg[31]~q ;
wire \phi_int_arr_reg[16]~q ;
wire \phi_int_arr_reg[17]~q ;
wire \phi_int_arr_reg[18]~q ;
wire \phi_int_arr_reg[19]~q ;
wire \phi_int_arr_reg[20]~q ;
wire \phi_int_arr_reg[21]~q ;
wire \phi_int_arr_reg[22]~q ;
wire \phi_int_arr_reg[23]~q ;
wire \phi_int_arr_reg[15]~q ;
wire \phi_int_arr_reg[14]~q ;
wire \phi_int_arr_reg[13]~q ;
wire \phi_int_arr_reg[12]~q ;
wire \phi_int_arr_reg[11]~q ;
wire \phi_int_arr_reg[10]~q ;
wire \phi_int_arr_reg[9]~q ;
wire \phi_int_arr_reg[8]~q ;
wire \phi_int_arr_reg[7]~q ;
wire \phi_int_arr_reg[6]~q ;
wire \phi_int_arr_reg[5]~q ;
wire \phi_int_arr_reg[4]~q ;
wire \phi_int_arr_reg[3]~q ;
wire \phi_int_arr_reg[2]~q ;
wire \phi_int_arr_reg[1]~q ;
wire \phi_int_arr_reg[0]~q ;


sine_lpm_add_sub_1 acc(
	.phi_int_arr_reg_24(\phi_int_arr_reg[24]~q ),
	.phi_int_arr_reg_25(\phi_int_arr_reg[25]~q ),
	.phi_int_arr_reg_26(\phi_int_arr_reg[26]~q ),
	.phi_int_arr_reg_27(\phi_int_arr_reg[27]~q ),
	.phi_int_arr_reg_28(\phi_int_arr_reg[28]~q ),
	.phi_int_arr_reg_29(\phi_int_arr_reg[29]~q ),
	.phi_int_arr_reg_30(\phi_int_arr_reg[30]~q ),
	.phi_int_arr_reg_31(\phi_int_arr_reg[31]~q ),
	.phi_int_arr_reg_16(\phi_int_arr_reg[16]~q ),
	.phi_int_arr_reg_17(\phi_int_arr_reg[17]~q ),
	.phi_int_arr_reg_18(\phi_int_arr_reg[18]~q ),
	.phi_int_arr_reg_19(\phi_int_arr_reg[19]~q ),
	.phi_int_arr_reg_20(\phi_int_arr_reg[20]~q ),
	.phi_int_arr_reg_21(\phi_int_arr_reg[21]~q ),
	.phi_int_arr_reg_22(\phi_int_arr_reg[22]~q ),
	.phi_int_arr_reg_23(\phi_int_arr_reg[23]~q ),
	.phi_int_arr_reg_15(\phi_int_arr_reg[15]~q ),
	.phi_int_arr_reg_14(\phi_int_arr_reg[14]~q ),
	.phi_int_arr_reg_13(\phi_int_arr_reg[13]~q ),
	.phi_int_arr_reg_12(\phi_int_arr_reg[12]~q ),
	.phi_int_arr_reg_11(\phi_int_arr_reg[11]~q ),
	.phi_int_arr_reg_10(\phi_int_arr_reg[10]~q ),
	.phi_int_arr_reg_9(\phi_int_arr_reg[9]~q ),
	.phi_int_arr_reg_8(\phi_int_arr_reg[8]~q ),
	.phi_int_arr_reg_7(\phi_int_arr_reg[7]~q ),
	.phi_int_arr_reg_6(\phi_int_arr_reg[6]~q ),
	.phi_int_arr_reg_5(\phi_int_arr_reg[5]~q ),
	.phi_int_arr_reg_4(\phi_int_arr_reg[4]~q ),
	.phi_int_arr_reg_3(\phi_int_arr_reg[3]~q ),
	.phi_int_arr_reg_2(\phi_int_arr_reg[2]~q ),
	.phi_int_arr_reg_1(\phi_int_arr_reg[1]~q ),
	.phi_int_arr_reg_0(\phi_int_arr_reg[0]~q ),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.clock(clk),
	.clken(clken),
	.reset_n(reset_n));

dffeas \phi_int_arr_reg[24] (
	.clk(clk),
	.d(pipeline_dffe_241),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[24]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[24] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[24] .power_up = "low";

dffeas \phi_int_arr_reg[25] (
	.clk(clk),
	.d(pipeline_dffe_251),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[25]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[25] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[25] .power_up = "low";

dffeas \phi_int_arr_reg[26] (
	.clk(clk),
	.d(pipeline_dffe_261),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[26]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[26] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[26] .power_up = "low";

dffeas \phi_int_arr_reg[27] (
	.clk(clk),
	.d(pipeline_dffe_271),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[27]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[27] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[27] .power_up = "low";

dffeas \phi_int_arr_reg[28] (
	.clk(clk),
	.d(pipeline_dffe_281),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[28]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[28] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[28] .power_up = "low";

dffeas \phi_int_arr_reg[29] (
	.clk(clk),
	.d(pipeline_dffe_291),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[29]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[29] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[29] .power_up = "low";

dffeas \phi_int_arr_reg[30] (
	.clk(clk),
	.d(pipeline_dffe_301),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[30]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[30] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[30] .power_up = "low";

dffeas \phi_int_arr_reg[31] (
	.clk(clk),
	.d(pipeline_dffe_311),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[31]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[31] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[31] .power_up = "low";

dffeas \phi_int_arr_reg[16] (
	.clk(clk),
	.d(pipeline_dffe_161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[16]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[16] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[16] .power_up = "low";

dffeas \phi_int_arr_reg[17] (
	.clk(clk),
	.d(pipeline_dffe_171),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[17]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[17] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[17] .power_up = "low";

dffeas \phi_int_arr_reg[18] (
	.clk(clk),
	.d(pipeline_dffe_181),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[18]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[18] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[18] .power_up = "low";

dffeas \phi_int_arr_reg[19] (
	.clk(clk),
	.d(pipeline_dffe_191),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[19]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[19] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[19] .power_up = "low";

dffeas \phi_int_arr_reg[20] (
	.clk(clk),
	.d(pipeline_dffe_201),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[20]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[20] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[20] .power_up = "low";

dffeas \phi_int_arr_reg[21] (
	.clk(clk),
	.d(pipeline_dffe_211),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[21]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[21] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[21] .power_up = "low";

dffeas \phi_int_arr_reg[22] (
	.clk(clk),
	.d(pipeline_dffe_221),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[22]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[22] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[22] .power_up = "low";

dffeas \phi_int_arr_reg[23] (
	.clk(clk),
	.d(pipeline_dffe_231),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[23]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[23] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[23] .power_up = "low";

dffeas \phi_int_arr_reg[15] (
	.clk(clk),
	.d(pipeline_dffe_151),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[15]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[15] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[15] .power_up = "low";

dffeas \phi_int_arr_reg[14] (
	.clk(clk),
	.d(pipeline_dffe_141),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[14]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[14] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[14] .power_up = "low";

dffeas \phi_int_arr_reg[13] (
	.clk(clk),
	.d(pipeline_dffe_131),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[13]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[13] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[13] .power_up = "low";

dffeas \phi_int_arr_reg[12] (
	.clk(clk),
	.d(pipeline_dffe_121),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[12]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[12] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[12] .power_up = "low";

dffeas \phi_int_arr_reg[11] (
	.clk(clk),
	.d(pipeline_dffe_111),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[11]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[11] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[11] .power_up = "low";

dffeas \phi_int_arr_reg[10] (
	.clk(clk),
	.d(pipeline_dffe_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[10]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[10] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[10] .power_up = "low";

dffeas \phi_int_arr_reg[9] (
	.clk(clk),
	.d(pipeline_dffe_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[9]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[9] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[9] .power_up = "low";

dffeas \phi_int_arr_reg[8] (
	.clk(clk),
	.d(pipeline_dffe_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[8]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[8] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[8] .power_up = "low";

dffeas \phi_int_arr_reg[7] (
	.clk(clk),
	.d(pipeline_dffe_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[7]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[7] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[7] .power_up = "low";

dffeas \phi_int_arr_reg[6] (
	.clk(clk),
	.d(pipeline_dffe_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[6]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[6] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[6] .power_up = "low";

dffeas \phi_int_arr_reg[5] (
	.clk(clk),
	.d(pipeline_dffe_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[5]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[5] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[5] .power_up = "low";

dffeas \phi_int_arr_reg[4] (
	.clk(clk),
	.d(pipeline_dffe_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[4]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[4] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[4] .power_up = "low";

dffeas \phi_int_arr_reg[3] (
	.clk(clk),
	.d(pipeline_dffe_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[3]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[3] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[3] .power_up = "low";

dffeas \phi_int_arr_reg[2] (
	.clk(clk),
	.d(pipeline_dffe_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[2]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[2] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[2] .power_up = "low";

dffeas \phi_int_arr_reg[1] (
	.clk(clk),
	.d(pipeline_dffe_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[1]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[1] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[1] .power_up = "low";

dffeas \phi_int_arr_reg[0] (
	.clk(clk),
	.d(pipeline_dffe_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_int_arr_reg[0]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[0] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[0] .power_up = "low";

endmodule

module sine_lpm_add_sub_1 (
	phi_int_arr_reg_24,
	phi_int_arr_reg_25,
	phi_int_arr_reg_26,
	phi_int_arr_reg_27,
	phi_int_arr_reg_28,
	phi_int_arr_reg_29,
	phi_int_arr_reg_30,
	phi_int_arr_reg_31,
	phi_int_arr_reg_16,
	phi_int_arr_reg_17,
	phi_int_arr_reg_18,
	phi_int_arr_reg_19,
	phi_int_arr_reg_20,
	phi_int_arr_reg_21,
	phi_int_arr_reg_22,
	phi_int_arr_reg_23,
	phi_int_arr_reg_15,
	phi_int_arr_reg_14,
	phi_int_arr_reg_13,
	phi_int_arr_reg_12,
	phi_int_arr_reg_11,
	phi_int_arr_reg_10,
	phi_int_arr_reg_9,
	phi_int_arr_reg_8,
	phi_int_arr_reg_7,
	phi_int_arr_reg_6,
	phi_int_arr_reg_5,
	phi_int_arr_reg_4,
	phi_int_arr_reg_3,
	phi_int_arr_reg_2,
	phi_int_arr_reg_1,
	phi_int_arr_reg_0,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	clock,
	clken,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	phi_int_arr_reg_24;
input 	phi_int_arr_reg_25;
input 	phi_int_arr_reg_26;
input 	phi_int_arr_reg_27;
input 	phi_int_arr_reg_28;
input 	phi_int_arr_reg_29;
input 	phi_int_arr_reg_30;
input 	phi_int_arr_reg_31;
input 	phi_int_arr_reg_16;
input 	phi_int_arr_reg_17;
input 	phi_int_arr_reg_18;
input 	phi_int_arr_reg_19;
input 	phi_int_arr_reg_20;
input 	phi_int_arr_reg_21;
input 	phi_int_arr_reg_22;
input 	phi_int_arr_reg_23;
input 	phi_int_arr_reg_15;
input 	phi_int_arr_reg_14;
input 	phi_int_arr_reg_13;
input 	phi_int_arr_reg_12;
input 	phi_int_arr_reg_11;
input 	phi_int_arr_reg_10;
input 	phi_int_arr_reg_9;
input 	phi_int_arr_reg_8;
input 	phi_int_arr_reg_7;
input 	phi_int_arr_reg_6;
input 	phi_int_arr_reg_5;
input 	phi_int_arr_reg_4;
input 	phi_int_arr_reg_3;
input 	phi_int_arr_reg_2;
input 	phi_int_arr_reg_1;
input 	phi_int_arr_reg_0;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
input 	clock;
input 	clken;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_add_sub_hth auto_generated(
	.phi_int_arr_reg_24(phi_int_arr_reg_24),
	.phi_int_arr_reg_25(phi_int_arr_reg_25),
	.phi_int_arr_reg_26(phi_int_arr_reg_26),
	.phi_int_arr_reg_27(phi_int_arr_reg_27),
	.phi_int_arr_reg_28(phi_int_arr_reg_28),
	.phi_int_arr_reg_29(phi_int_arr_reg_29),
	.phi_int_arr_reg_30(phi_int_arr_reg_30),
	.phi_int_arr_reg_31(phi_int_arr_reg_31),
	.phi_int_arr_reg_16(phi_int_arr_reg_16),
	.phi_int_arr_reg_17(phi_int_arr_reg_17),
	.phi_int_arr_reg_18(phi_int_arr_reg_18),
	.phi_int_arr_reg_19(phi_int_arr_reg_19),
	.phi_int_arr_reg_20(phi_int_arr_reg_20),
	.phi_int_arr_reg_21(phi_int_arr_reg_21),
	.phi_int_arr_reg_22(phi_int_arr_reg_22),
	.phi_int_arr_reg_23(phi_int_arr_reg_23),
	.phi_int_arr_reg_15(phi_int_arr_reg_15),
	.phi_int_arr_reg_14(phi_int_arr_reg_14),
	.phi_int_arr_reg_13(phi_int_arr_reg_13),
	.phi_int_arr_reg_12(phi_int_arr_reg_12),
	.phi_int_arr_reg_11(phi_int_arr_reg_11),
	.phi_int_arr_reg_10(phi_int_arr_reg_10),
	.phi_int_arr_reg_9(phi_int_arr_reg_9),
	.phi_int_arr_reg_8(phi_int_arr_reg_8),
	.phi_int_arr_reg_7(phi_int_arr_reg_7),
	.phi_int_arr_reg_6(phi_int_arr_reg_6),
	.phi_int_arr_reg_5(phi_int_arr_reg_5),
	.phi_int_arr_reg_4(phi_int_arr_reg_4),
	.phi_int_arr_reg_3(phi_int_arr_reg_3),
	.phi_int_arr_reg_2(phi_int_arr_reg_2),
	.phi_int_arr_reg_1(phi_int_arr_reg_1),
	.phi_int_arr_reg_0(phi_int_arr_reg_0),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.clock(clock),
	.clken(clken),
	.reset_n(reset_n));

endmodule

module sine_add_sub_hth (
	phi_int_arr_reg_24,
	phi_int_arr_reg_25,
	phi_int_arr_reg_26,
	phi_int_arr_reg_27,
	phi_int_arr_reg_28,
	phi_int_arr_reg_29,
	phi_int_arr_reg_30,
	phi_int_arr_reg_31,
	phi_int_arr_reg_16,
	phi_int_arr_reg_17,
	phi_int_arr_reg_18,
	phi_int_arr_reg_19,
	phi_int_arr_reg_20,
	phi_int_arr_reg_21,
	phi_int_arr_reg_22,
	phi_int_arr_reg_23,
	phi_int_arr_reg_15,
	phi_int_arr_reg_14,
	phi_int_arr_reg_13,
	phi_int_arr_reg_12,
	phi_int_arr_reg_11,
	phi_int_arr_reg_10,
	phi_int_arr_reg_9,
	phi_int_arr_reg_8,
	phi_int_arr_reg_7,
	phi_int_arr_reg_6,
	phi_int_arr_reg_5,
	phi_int_arr_reg_4,
	phi_int_arr_reg_3,
	phi_int_arr_reg_2,
	phi_int_arr_reg_1,
	phi_int_arr_reg_0,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	clock,
	clken,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	phi_int_arr_reg_24;
input 	phi_int_arr_reg_25;
input 	phi_int_arr_reg_26;
input 	phi_int_arr_reg_27;
input 	phi_int_arr_reg_28;
input 	phi_int_arr_reg_29;
input 	phi_int_arr_reg_30;
input 	phi_int_arr_reg_31;
input 	phi_int_arr_reg_16;
input 	phi_int_arr_reg_17;
input 	phi_int_arr_reg_18;
input 	phi_int_arr_reg_19;
input 	phi_int_arr_reg_20;
input 	phi_int_arr_reg_21;
input 	phi_int_arr_reg_22;
input 	phi_int_arr_reg_23;
input 	phi_int_arr_reg_15;
input 	phi_int_arr_reg_14;
input 	phi_int_arr_reg_13;
input 	phi_int_arr_reg_12;
input 	phi_int_arr_reg_11;
input 	phi_int_arr_reg_10;
input 	phi_int_arr_reg_9;
input 	phi_int_arr_reg_8;
input 	phi_int_arr_reg_7;
input 	phi_int_arr_reg_6;
input 	phi_int_arr_reg_5;
input 	phi_int_arr_reg_4;
input 	phi_int_arr_reg_3;
input 	phi_int_arr_reg_2;
input 	phi_int_arr_reg_1;
input 	phi_int_arr_reg_0;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
input 	clock;
input 	clken;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~125_sumout ;
wire \pipeline_dffe[0]~q ;
wire \op_1~126 ;
wire \op_1~121_sumout ;
wire \pipeline_dffe[1]~q ;
wire \op_1~122 ;
wire \op_1~117_sumout ;
wire \pipeline_dffe[2]~q ;
wire \op_1~118 ;
wire \op_1~113_sumout ;
wire \pipeline_dffe[3]~q ;
wire \op_1~114 ;
wire \op_1~109_sumout ;
wire \pipeline_dffe[4]~q ;
wire \op_1~110 ;
wire \op_1~105_sumout ;
wire \pipeline_dffe[5]~q ;
wire \op_1~106 ;
wire \op_1~101_sumout ;
wire \pipeline_dffe[6]~q ;
wire \op_1~102 ;
wire \op_1~97_sumout ;
wire \pipeline_dffe[7]~q ;
wire \op_1~98 ;
wire \op_1~93_sumout ;
wire \pipeline_dffe[8]~q ;
wire \op_1~94 ;
wire \op_1~89_sumout ;
wire \pipeline_dffe[9]~q ;
wire \op_1~90 ;
wire \op_1~85_sumout ;
wire \pipeline_dffe[10]~q ;
wire \op_1~86 ;
wire \op_1~82 ;
wire \op_1~78 ;
wire \op_1~74 ;
wire \op_1~70 ;
wire \op_1~66 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~50 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~6 ;
wire \op_1~9_sumout ;
wire \op_1~10 ;
wire \op_1~13_sumout ;
wire \op_1~14 ;
wire \op_1~17_sumout ;
wire \op_1~18 ;
wire \op_1~21_sumout ;
wire \op_1~22 ;
wire \op_1~25_sumout ;
wire \op_1~26 ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~73_sumout ;
wire \op_1~77_sumout ;
wire \op_1~81_sumout ;


dffeas \pipeline_dffe[24] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_24),
	.prn(vcc));
defparam \pipeline_dffe[24] .is_wysiwyg = "true";
defparam \pipeline_dffe[24] .power_up = "low";

dffeas \pipeline_dffe[25] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_25),
	.prn(vcc));
defparam \pipeline_dffe[25] .is_wysiwyg = "true";
defparam \pipeline_dffe[25] .power_up = "low";

dffeas \pipeline_dffe[26] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_26),
	.prn(vcc));
defparam \pipeline_dffe[26] .is_wysiwyg = "true";
defparam \pipeline_dffe[26] .power_up = "low";

dffeas \pipeline_dffe[27] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_27),
	.prn(vcc));
defparam \pipeline_dffe[27] .is_wysiwyg = "true";
defparam \pipeline_dffe[27] .power_up = "low";

dffeas \pipeline_dffe[28] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_28),
	.prn(vcc));
defparam \pipeline_dffe[28] .is_wysiwyg = "true";
defparam \pipeline_dffe[28] .power_up = "low";

dffeas \pipeline_dffe[29] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_29),
	.prn(vcc));
defparam \pipeline_dffe[29] .is_wysiwyg = "true";
defparam \pipeline_dffe[29] .power_up = "low";

dffeas \pipeline_dffe[30] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_30),
	.prn(vcc));
defparam \pipeline_dffe[30] .is_wysiwyg = "true";
defparam \pipeline_dffe[30] .power_up = "low";

dffeas \pipeline_dffe[31] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_31),
	.prn(vcc));
defparam \pipeline_dffe[31] .is_wysiwyg = "true";
defparam \pipeline_dffe[31] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[18] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \pipeline_dffe[18] .is_wysiwyg = "true";
defparam \pipeline_dffe[18] .power_up = "low";

dffeas \pipeline_dffe[19] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \pipeline_dffe[19] .is_wysiwyg = "true";
defparam \pipeline_dffe[19] .power_up = "low";

dffeas \pipeline_dffe[20] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_20),
	.prn(vcc));
defparam \pipeline_dffe[20] .is_wysiwyg = "true";
defparam \pipeline_dffe[20] .power_up = "low";

dffeas \pipeline_dffe[21] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_21),
	.prn(vcc));
defparam \pipeline_dffe[21] .is_wysiwyg = "true";
defparam \pipeline_dffe[21] .power_up = "low";

dffeas \pipeline_dffe[22] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_22),
	.prn(vcc));
defparam \pipeline_dffe[22] .is_wysiwyg = "true";
defparam \pipeline_dffe[22] .power_up = "low";

dffeas \pipeline_dffe[23] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_23),
	.prn(vcc));
defparam \pipeline_dffe[23] .is_wysiwyg = "true";
defparam \pipeline_dffe[23] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~73_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~77_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~81_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

cyclonev_lcell_comb \op_1~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_0),
	.datae(gnd),
	.dataf(!\pipeline_dffe[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~125_sumout ),
	.cout(\op_1~126 ),
	.shareout());
defparam \op_1~125 .extended_lut = "off";
defparam \op_1~125 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~125 .shared_arith = "off";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~125_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[0]~q ),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

cyclonev_lcell_comb \op_1~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_1),
	.datae(gnd),
	.dataf(!\pipeline_dffe[1]~q ),
	.datag(gnd),
	.cin(\op_1~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~121_sumout ),
	.cout(\op_1~122 ),
	.shareout());
defparam \op_1~121 .extended_lut = "off";
defparam \op_1~121 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~121 .shared_arith = "off";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~121_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[1]~q ),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

cyclonev_lcell_comb \op_1~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_2),
	.datae(gnd),
	.dataf(!\pipeline_dffe[2]~q ),
	.datag(gnd),
	.cin(\op_1~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~117_sumout ),
	.cout(\op_1~118 ),
	.shareout());
defparam \op_1~117 .extended_lut = "off";
defparam \op_1~117 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~117 .shared_arith = "off";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~117_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[2]~q ),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

cyclonev_lcell_comb \op_1~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_3),
	.datae(gnd),
	.dataf(!\pipeline_dffe[3]~q ),
	.datag(gnd),
	.cin(\op_1~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~113_sumout ),
	.cout(\op_1~114 ),
	.shareout());
defparam \op_1~113 .extended_lut = "off";
defparam \op_1~113 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~113 .shared_arith = "off";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~113_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[3]~q ),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

cyclonev_lcell_comb \op_1~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_4),
	.datae(gnd),
	.dataf(!\pipeline_dffe[4]~q ),
	.datag(gnd),
	.cin(\op_1~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~109_sumout ),
	.cout(\op_1~110 ),
	.shareout());
defparam \op_1~109 .extended_lut = "off";
defparam \op_1~109 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~109 .shared_arith = "off";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~109_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[4]~q ),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

cyclonev_lcell_comb \op_1~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_5),
	.datae(gnd),
	.dataf(!\pipeline_dffe[5]~q ),
	.datag(gnd),
	.cin(\op_1~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~105_sumout ),
	.cout(\op_1~106 ),
	.shareout());
defparam \op_1~105 .extended_lut = "off";
defparam \op_1~105 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~105 .shared_arith = "off";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~105_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[5]~q ),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

cyclonev_lcell_comb \op_1~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_6),
	.datae(gnd),
	.dataf(!\pipeline_dffe[6]~q ),
	.datag(gnd),
	.cin(\op_1~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~101_sumout ),
	.cout(\op_1~102 ),
	.shareout());
defparam \op_1~101 .extended_lut = "off";
defparam \op_1~101 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~101 .shared_arith = "off";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~101_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[6]~q ),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

cyclonev_lcell_comb \op_1~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_7),
	.datae(gnd),
	.dataf(!\pipeline_dffe[7]~q ),
	.datag(gnd),
	.cin(\op_1~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~97_sumout ),
	.cout(\op_1~98 ),
	.shareout());
defparam \op_1~97 .extended_lut = "off";
defparam \op_1~97 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~97 .shared_arith = "off";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~97_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[7]~q ),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

cyclonev_lcell_comb \op_1~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_8),
	.datae(gnd),
	.dataf(!\pipeline_dffe[8]~q ),
	.datag(gnd),
	.cin(\op_1~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~93_sumout ),
	.cout(\op_1~94 ),
	.shareout());
defparam \op_1~93 .extended_lut = "off";
defparam \op_1~93 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~93 .shared_arith = "off";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~93_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[8]~q ),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

cyclonev_lcell_comb \op_1~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_9),
	.datae(gnd),
	.dataf(!\pipeline_dffe[9]~q ),
	.datag(gnd),
	.cin(\op_1~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~89_sumout ),
	.cout(\op_1~90 ),
	.shareout());
defparam \op_1~89 .extended_lut = "off";
defparam \op_1~89 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~89 .shared_arith = "off";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~89_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[9]~q ),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

cyclonev_lcell_comb \op_1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_10),
	.datae(gnd),
	.dataf(!\pipeline_dffe[10]~q ),
	.datag(gnd),
	.cin(\op_1~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~85_sumout ),
	.cout(\op_1~86 ),
	.shareout());
defparam \op_1~85 .extended_lut = "off";
defparam \op_1~85 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~85 .shared_arith = "off";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~85_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[10]~q ),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

cyclonev_lcell_comb \op_1~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_11),
	.datae(gnd),
	.dataf(!pipeline_dffe_11),
	.datag(gnd),
	.cin(\op_1~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~81_sumout ),
	.cout(\op_1~82 ),
	.shareout());
defparam \op_1~81 .extended_lut = "off";
defparam \op_1~81 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~81 .shared_arith = "off";

cyclonev_lcell_comb \op_1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_12),
	.datae(gnd),
	.dataf(!pipeline_dffe_12),
	.datag(gnd),
	.cin(\op_1~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~77_sumout ),
	.cout(\op_1~78 ),
	.shareout());
defparam \op_1~77 .extended_lut = "off";
defparam \op_1~77 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~77 .shared_arith = "off";

cyclonev_lcell_comb \op_1~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_13),
	.datae(gnd),
	.dataf(!pipeline_dffe_13),
	.datag(gnd),
	.cin(\op_1~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~73_sumout ),
	.cout(\op_1~74 ),
	.shareout());
defparam \op_1~73 .extended_lut = "off";
defparam \op_1~73 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~73 .shared_arith = "off";

cyclonev_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_14),
	.datae(gnd),
	.dataf(!pipeline_dffe_14),
	.datag(gnd),
	.cin(\op_1~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

cyclonev_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_15),
	.datae(gnd),
	.dataf(!pipeline_dffe_15),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_16),
	.datae(gnd),
	.dataf(!pipeline_dffe_16),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_17),
	.datae(gnd),
	.dataf(!pipeline_dffe_17),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_18),
	.datae(gnd),
	.dataf(!pipeline_dffe_18),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_19),
	.datae(gnd),
	.dataf(!pipeline_dffe_19),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_20),
	.datae(gnd),
	.dataf(!pipeline_dffe_20),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

cyclonev_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_21),
	.datae(gnd),
	.dataf(!pipeline_dffe_21),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

cyclonev_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_22),
	.datae(gnd),
	.dataf(!pipeline_dffe_22),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

cyclonev_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_23),
	.datae(gnd),
	.dataf(!pipeline_dffe_23),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_24),
	.datae(gnd),
	.dataf(!pipeline_dffe_24),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_25),
	.datae(gnd),
	.dataf(!pipeline_dffe_25),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_26),
	.datae(gnd),
	.dataf(!pipeline_dffe_26),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_27),
	.datae(gnd),
	.dataf(!pipeline_dffe_27),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_28),
	.datae(gnd),
	.dataf(!pipeline_dffe_28),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_29),
	.datae(gnd),
	.dataf(!pipeline_dffe_29),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_30),
	.datae(gnd),
	.dataf(!pipeline_dffe_30),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_31),
	.datae(gnd),
	.dataf(!pipeline_dffe_31),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

endmodule

module sine_asj_dxx (
	dxxpdo_13,
	dxxpdo_14,
	dxxpdo_15,
	dxxpdo_16,
	dxxpdo_17,
	dxxpdo_18,
	dxxpdo_19,
	dxxpdo_20,
	dxxpdo_5,
	dxxpdo_6,
	dxxpdo_7,
	dxxpdo_8,
	dxxpdo_9,
	dxxpdo_10,
	dxxpdo_11,
	dxxpdo_12,
	dxxrv_3,
	dxxrv_2,
	dxxrv_1,
	dxxrv_0,
	result_a_28,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	NJQG9082,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dxxpdo_13;
output 	dxxpdo_14;
output 	dxxpdo_15;
output 	dxxpdo_16;
output 	dxxpdo_17;
output 	dxxpdo_18;
output 	dxxpdo_19;
output 	dxxpdo_20;
output 	dxxpdo_5;
output 	dxxpdo_6;
output 	dxxpdo_7;
output 	dxxpdo_8;
output 	dxxpdo_9;
output 	dxxpdo_10;
output 	dxxpdo_11;
output 	dxxpdo_12;
input 	dxxrv_3;
input 	dxxrv_2;
input 	dxxrv_1;
input 	dxxrv_0;
input 	result_a_28;
input 	pipeline_dffe_24;
input 	pipeline_dffe_25;
input 	pipeline_dffe_26;
input 	pipeline_dffe_27;
input 	pipeline_dffe_28;
input 	pipeline_dffe_29;
input 	pipeline_dffe_30;
input 	pipeline_dffe_31;
input 	pipeline_dffe_16;
input 	pipeline_dffe_17;
input 	pipeline_dffe_18;
input 	pipeline_dffe_19;
input 	pipeline_dffe_20;
input 	pipeline_dffe_21;
input 	pipeline_dffe_22;
input 	pipeline_dffe_23;
input 	pipeline_dffe_15;
input 	pipeline_dffe_14;
input 	pipeline_dffe_13;
input 	pipeline_dffe_12;
input 	pipeline_dffe_11;
input 	NJQG9082;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~82_cout ;
wire \Add0~78_cout ;
wire \Add0~74_cout ;
wire \Add0~70_cout ;
wire \Add0~66_cout ;
wire \Add0~34 ;
wire \Add0~38 ;
wire \Add0~42 ;
wire \Add0~46 ;
wire \Add0~50 ;
wire \Add0~54 ;
wire \Add0~58 ;
wire \Add0~62 ;
wire \Add0~1_sumout ;
wire \phi_dither_out_w[13]~q ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \phi_dither_out_w[14]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \phi_dither_out_w[15]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \phi_dither_out_w[16]~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \phi_dither_out_w[17]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \phi_dither_out_w[18]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \phi_dither_out_w[19]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \phi_dither_out_w[20]~q ;
wire \Add0~33_sumout ;
wire \phi_dither_out_w[5]~q ;
wire \Add0~37_sumout ;
wire \phi_dither_out_w[6]~q ;
wire \Add0~41_sumout ;
wire \phi_dither_out_w[7]~q ;
wire \Add0~45_sumout ;
wire \phi_dither_out_w[8]~q ;
wire \Add0~49_sumout ;
wire \phi_dither_out_w[9]~q ;
wire \Add0~53_sumout ;
wire \phi_dither_out_w[10]~q ;
wire \Add0~57_sumout ;
wire \phi_dither_out_w[11]~q ;
wire \Add0~61_sumout ;
wire \phi_dither_out_w[12]~q ;


dffeas \dxxpdo[13] (
	.clk(clk),
	.d(\phi_dither_out_w[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_13),
	.prn(vcc));
defparam \dxxpdo[13] .is_wysiwyg = "true";
defparam \dxxpdo[13] .power_up = "low";

dffeas \dxxpdo[14] (
	.clk(clk),
	.d(\phi_dither_out_w[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_14),
	.prn(vcc));
defparam \dxxpdo[14] .is_wysiwyg = "true";
defparam \dxxpdo[14] .power_up = "low";

dffeas \dxxpdo[15] (
	.clk(clk),
	.d(\phi_dither_out_w[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_15),
	.prn(vcc));
defparam \dxxpdo[15] .is_wysiwyg = "true";
defparam \dxxpdo[15] .power_up = "low";

dffeas \dxxpdo[16] (
	.clk(clk),
	.d(\phi_dither_out_w[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_16),
	.prn(vcc));
defparam \dxxpdo[16] .is_wysiwyg = "true";
defparam \dxxpdo[16] .power_up = "low";

dffeas \dxxpdo[17] (
	.clk(clk),
	.d(\phi_dither_out_w[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_17),
	.prn(vcc));
defparam \dxxpdo[17] .is_wysiwyg = "true";
defparam \dxxpdo[17] .power_up = "low";

dffeas \dxxpdo[18] (
	.clk(clk),
	.d(\phi_dither_out_w[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_18),
	.prn(vcc));
defparam \dxxpdo[18] .is_wysiwyg = "true";
defparam \dxxpdo[18] .power_up = "low";

dffeas \dxxpdo[19] (
	.clk(clk),
	.d(\phi_dither_out_w[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_19),
	.prn(vcc));
defparam \dxxpdo[19] .is_wysiwyg = "true";
defparam \dxxpdo[19] .power_up = "low";

dffeas \dxxpdo[20] (
	.clk(clk),
	.d(\phi_dither_out_w[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_20),
	.prn(vcc));
defparam \dxxpdo[20] .is_wysiwyg = "true";
defparam \dxxpdo[20] .power_up = "low";

dffeas \dxxpdo[5] (
	.clk(clk),
	.d(\phi_dither_out_w[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_5),
	.prn(vcc));
defparam \dxxpdo[5] .is_wysiwyg = "true";
defparam \dxxpdo[5] .power_up = "low";

dffeas \dxxpdo[6] (
	.clk(clk),
	.d(\phi_dither_out_w[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_6),
	.prn(vcc));
defparam \dxxpdo[6] .is_wysiwyg = "true";
defparam \dxxpdo[6] .power_up = "low";

dffeas \dxxpdo[7] (
	.clk(clk),
	.d(\phi_dither_out_w[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_7),
	.prn(vcc));
defparam \dxxpdo[7] .is_wysiwyg = "true";
defparam \dxxpdo[7] .power_up = "low";

dffeas \dxxpdo[8] (
	.clk(clk),
	.d(\phi_dither_out_w[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_8),
	.prn(vcc));
defparam \dxxpdo[8] .is_wysiwyg = "true";
defparam \dxxpdo[8] .power_up = "low";

dffeas \dxxpdo[9] (
	.clk(clk),
	.d(\phi_dither_out_w[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_9),
	.prn(vcc));
defparam \dxxpdo[9] .is_wysiwyg = "true";
defparam \dxxpdo[9] .power_up = "low";

dffeas \dxxpdo[10] (
	.clk(clk),
	.d(\phi_dither_out_w[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_10),
	.prn(vcc));
defparam \dxxpdo[10] .is_wysiwyg = "true";
defparam \dxxpdo[10] .power_up = "low";

dffeas \dxxpdo[11] (
	.clk(clk),
	.d(\phi_dither_out_w[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_11),
	.prn(vcc));
defparam \dxxpdo[11] .is_wysiwyg = "true";
defparam \dxxpdo[11] .power_up = "low";

dffeas \dxxpdo[12] (
	.clk(clk),
	.d(\phi_dither_out_w[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxpdo_12),
	.prn(vcc));
defparam \dxxpdo[12] .is_wysiwyg = "true";
defparam \dxxpdo[12] .power_up = "low";

cyclonev_lcell_comb \Add0~82 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_0),
	.datae(gnd),
	.dataf(!pipeline_dffe_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~82_cout ),
	.shareout());
defparam \Add0~82 .extended_lut = "off";
defparam \Add0~82 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~82 .shared_arith = "off";

cyclonev_lcell_comb \Add0~78 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_1),
	.datae(gnd),
	.dataf(!pipeline_dffe_12),
	.datag(gnd),
	.cin(\Add0~82_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~78_cout ),
	.shareout());
defparam \Add0~78 .extended_lut = "off";
defparam \Add0~78 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~78 .shared_arith = "off";

cyclonev_lcell_comb \Add0~74 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_2),
	.datae(gnd),
	.dataf(!pipeline_dffe_13),
	.datag(gnd),
	.cin(\Add0~78_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~74_cout ),
	.shareout());
defparam \Add0~74 .extended_lut = "off";
defparam \Add0~74 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~74 .shared_arith = "off";

cyclonev_lcell_comb \Add0~70 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_14),
	.datag(gnd),
	.cin(\Add0~74_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~70_cout ),
	.shareout());
defparam \Add0~70 .extended_lut = "off";
defparam \Add0~70 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~70 .shared_arith = "off";

cyclonev_lcell_comb \Add0~66 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_15),
	.datag(gnd),
	.cin(\Add0~70_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~66_cout ),
	.shareout());
defparam \Add0~66 .extended_lut = "off";
defparam \Add0~66 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~66 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_16),
	.datag(gnd),
	.cin(\Add0~66_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_17),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_18),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_19),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~45 .shared_arith = "off";

cyclonev_lcell_comb \Add0~49 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_20),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~49 .shared_arith = "off";

cyclonev_lcell_comb \Add0~53 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_21),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~53 .shared_arith = "off";

cyclonev_lcell_comb \Add0~57 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_22),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~57 .shared_arith = "off";

cyclonev_lcell_comb \Add0~61 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_23),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~61 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_24),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \phi_dither_out_w[13] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[13]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[13] .is_wysiwyg = "true";
defparam \phi_dither_out_w[13] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_25),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \phi_dither_out_w[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[14]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[14] .is_wysiwyg = "true";
defparam \phi_dither_out_w[14] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_26),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \phi_dither_out_w[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[15]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[15] .is_wysiwyg = "true";
defparam \phi_dither_out_w[15] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_27),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \phi_dither_out_w[16] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[16]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[16] .is_wysiwyg = "true";
defparam \phi_dither_out_w[16] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_28),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \phi_dither_out_w[17] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[17]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[17] .is_wysiwyg = "true";
defparam \phi_dither_out_w[17] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_29),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \phi_dither_out_w[18] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[18]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[18] .is_wysiwyg = "true";
defparam \phi_dither_out_w[18] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_30),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \phi_dither_out_w[19] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[19]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[19] .is_wysiwyg = "true";
defparam \phi_dither_out_w[19] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_31),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \phi_dither_out_w[20] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[20]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[20] .is_wysiwyg = "true";
defparam \phi_dither_out_w[20] .power_up = "low";

dffeas \phi_dither_out_w[5] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[5]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[5] .is_wysiwyg = "true";
defparam \phi_dither_out_w[5] .power_up = "low";

dffeas \phi_dither_out_w[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[6]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[6] .is_wysiwyg = "true";
defparam \phi_dither_out_w[6] .power_up = "low";

dffeas \phi_dither_out_w[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[7]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[7] .is_wysiwyg = "true";
defparam \phi_dither_out_w[7] .power_up = "low";

dffeas \phi_dither_out_w[8] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[8]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[8] .is_wysiwyg = "true";
defparam \phi_dither_out_w[8] .power_up = "low";

dffeas \phi_dither_out_w[9] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[9]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[9] .is_wysiwyg = "true";
defparam \phi_dither_out_w[9] .power_up = "low";

dffeas \phi_dither_out_w[10] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[10]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[10] .is_wysiwyg = "true";
defparam \phi_dither_out_w[10] .power_up = "low";

dffeas \phi_dither_out_w[11] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[11]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[11] .is_wysiwyg = "true";
defparam \phi_dither_out_w[11] .power_up = "low";

dffeas \phi_dither_out_w[12] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_dither_out_w[12]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[12] .is_wysiwyg = "true";
defparam \phi_dither_out_w[12] .power_up = "low";

endmodule

module sine_asj_dxx_g (
	dxxrv_3,
	dxxrv_2,
	dxxrv_1,
	dxxrv_0,
	result_a_28,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dxxrv_3;
output 	dxxrv_2;
output 	dxxrv_1;
output 	dxxrv_0;
input 	result_a_28;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lsfr_reg~10_combout ;
wire \lsfr_reg[0]~q ;
wire \lsfr_reg[1]~q ;
wire \lsfr_reg~9_combout ;
wire \lsfr_reg[2]~q ;
wire \lsfr_reg~8_combout ;
wire \lsfr_reg[3]~q ;
wire \lsfr_reg~7_combout ;
wire \lsfr_reg[4]~q ;
wire \lsfr_reg[5]~q ;
wire \lsfr_reg~6_combout ;
wire \lsfr_reg[6]~q ;
wire \lsfr_reg~5_combout ;
wire \lsfr_reg[7]~q ;
wire \lsfr_reg[8]~q ;
wire \lsfr_reg~3_combout ;
wire \lsfr_reg[9]~q ;
wire \lsfr_reg[10]~q ;
wire \lsfr_reg~2_combout ;
wire \lsfr_reg[11]~q ;
wire \lsfr_reg~1_combout ;
wire \lsfr_reg[12]~q ;
wire \lsfr_reg[13]~q ;
wire \lsfr_reg[14]~q ;
wire \lsfr_reg~0_combout ;
wire \lsfr_reg[15]~q ;
wire \Add0~0_combout ;
wire \Add0~1_combout ;
wire \Add0~2_combout ;
wire \lsfr_reg~4_combout ;


dffeas \dxxrv[3] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxrv_3),
	.prn(vcc));
defparam \dxxrv[3] .is_wysiwyg = "true";
defparam \dxxrv[3] .power_up = "low";

dffeas \dxxrv[2] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxrv_2),
	.prn(vcc));
defparam \dxxrv[2] .is_wysiwyg = "true";
defparam \dxxrv[2] .power_up = "low";

dffeas \dxxrv[1] (
	.clk(clk),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxrv_1),
	.prn(vcc));
defparam \dxxrv[1] .is_wysiwyg = "true";
defparam \dxxrv[1] .power_up = "low";

dffeas \dxxrv[0] (
	.clk(clk),
	.d(\lsfr_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(dxxrv_0),
	.prn(vcc));
defparam \dxxrv[0] .is_wysiwyg = "true";
defparam \dxxrv[0] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~10 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[14]~q ),
	.datac(!\lsfr_reg[12]~q ),
	.datad(!\lsfr_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~10 .extended_lut = "off";
defparam \lsfr_reg~10 .lut_mask = 64'h6996699669966996;
defparam \lsfr_reg~10 .shared_arith = "off";

dffeas \lsfr_reg[0] (
	.clk(clk),
	.d(\lsfr_reg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(result_a_28),
	.q(\lsfr_reg[0]~q ),
	.prn(vcc));
defparam \lsfr_reg[0] .is_wysiwyg = "true";
defparam \lsfr_reg[0] .power_up = "low";

dffeas \lsfr_reg[1] (
	.clk(clk),
	.d(\lsfr_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[1]~q ),
	.prn(vcc));
defparam \lsfr_reg[1] .is_wysiwyg = "true";
defparam \lsfr_reg[1] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~9 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~9 .extended_lut = "off";
defparam \lsfr_reg~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~9 .shared_arith = "off";

dffeas \lsfr_reg[2] (
	.clk(clk),
	.d(\lsfr_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[2]~q ),
	.prn(vcc));
defparam \lsfr_reg[2] .is_wysiwyg = "true";
defparam \lsfr_reg[2] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~8 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~8 .extended_lut = "off";
defparam \lsfr_reg~8 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~8 .shared_arith = "off";

dffeas \lsfr_reg[3] (
	.clk(clk),
	.d(\lsfr_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[3]~q ),
	.prn(vcc));
defparam \lsfr_reg[3] .is_wysiwyg = "true";
defparam \lsfr_reg[3] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~7 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~7 .extended_lut = "off";
defparam \lsfr_reg~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~7 .shared_arith = "off";

dffeas \lsfr_reg[4] (
	.clk(clk),
	.d(\lsfr_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[4]~q ),
	.prn(vcc));
defparam \lsfr_reg[4] .is_wysiwyg = "true";
defparam \lsfr_reg[4] .power_up = "low";

dffeas \lsfr_reg[5] (
	.clk(clk),
	.d(\lsfr_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[5]~q ),
	.prn(vcc));
defparam \lsfr_reg[5] .is_wysiwyg = "true";
defparam \lsfr_reg[5] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~6 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~6 .extended_lut = "off";
defparam \lsfr_reg~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~6 .shared_arith = "off";

dffeas \lsfr_reg[6] (
	.clk(clk),
	.d(\lsfr_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[6]~q ),
	.prn(vcc));
defparam \lsfr_reg[6] .is_wysiwyg = "true";
defparam \lsfr_reg[6] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~5 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~5 .extended_lut = "off";
defparam \lsfr_reg~5 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~5 .shared_arith = "off";

dffeas \lsfr_reg[7] (
	.clk(clk),
	.d(\lsfr_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[7]~q ),
	.prn(vcc));
defparam \lsfr_reg[7] .is_wysiwyg = "true";
defparam \lsfr_reg[7] .power_up = "low";

dffeas \lsfr_reg[8] (
	.clk(clk),
	.d(\lsfr_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[8]~q ),
	.prn(vcc));
defparam \lsfr_reg[8] .is_wysiwyg = "true";
defparam \lsfr_reg[8] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~3 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~3 .extended_lut = "off";
defparam \lsfr_reg~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~3 .shared_arith = "off";

dffeas \lsfr_reg[9] (
	.clk(clk),
	.d(\lsfr_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[9]~q ),
	.prn(vcc));
defparam \lsfr_reg[9] .is_wysiwyg = "true";
defparam \lsfr_reg[9] .power_up = "low";

dffeas \lsfr_reg[10] (
	.clk(clk),
	.d(\lsfr_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[10]~q ),
	.prn(vcc));
defparam \lsfr_reg[10] .is_wysiwyg = "true";
defparam \lsfr_reg[10] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~2 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~2 .extended_lut = "off";
defparam \lsfr_reg~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~2 .shared_arith = "off";

dffeas \lsfr_reg[11] (
	.clk(clk),
	.d(\lsfr_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[11]~q ),
	.prn(vcc));
defparam \lsfr_reg[11] .is_wysiwyg = "true";
defparam \lsfr_reg[11] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~1 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~1 .extended_lut = "off";
defparam \lsfr_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~1 .shared_arith = "off";

dffeas \lsfr_reg[12] (
	.clk(clk),
	.d(\lsfr_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[12]~q ),
	.prn(vcc));
defparam \lsfr_reg[12] .is_wysiwyg = "true";
defparam \lsfr_reg[12] .power_up = "low";

dffeas \lsfr_reg[13] (
	.clk(clk),
	.d(\lsfr_reg[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[13]~q ),
	.prn(vcc));
defparam \lsfr_reg[13] .is_wysiwyg = "true";
defparam \lsfr_reg[13] .power_up = "low";

dffeas \lsfr_reg[14] (
	.clk(clk),
	.d(\lsfr_reg[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[14]~q ),
	.prn(vcc));
defparam \lsfr_reg[14] .is_wysiwyg = "true";
defparam \lsfr_reg[14] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~0 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~0 .extended_lut = "off";
defparam \lsfr_reg~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~0 .shared_arith = "off";

dffeas \lsfr_reg[15] (
	.clk(clk),
	.d(\lsfr_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(result_a_28),
	.q(\lsfr_reg[15]~q ),
	.prn(vcc));
defparam \lsfr_reg[15] .is_wysiwyg = "true";
defparam \lsfr_reg[15] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[14]~q ),
	.datac(!\lsfr_reg[13]~q ),
	.datad(!\lsfr_reg[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[14]~q ),
	.datac(!\lsfr_reg[13]~q ),
	.datad(!\lsfr_reg[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6996699669966996;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[13]~q ),
	.datac(!\lsfr_reg[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h9696969696969696;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \lsfr_reg~4 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~4 .extended_lut = "off";
defparam \lsfr_reg~4 .lut_mask = 64'h6666666666666666;
defparam \lsfr_reg~4 .shared_arith = "off";

endmodule

module sine_asj_gam_dp (
	rom_add_cc_temp_0,
	rom_add_cc_temp_1,
	rom_add_cc_temp_2,
	rom_add_cc_temp_3,
	rom_add_cc_temp_4,
	rom_add_cc_temp_5,
	rom_add_cs_6,
	rom_add_cs_7,
	rom_add_cc_temp_6,
	rom_add_cc_temp_7,
	rom_add_f_0,
	rom_add_f_1,
	rom_add_f_2,
	rom_add_f_3,
	rom_add_f_4,
	rom_add_f_5,
	rom_add_f_6,
	rom_add_f_7,
	result_a_28,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	rom_add_cc_temp_0;
output 	rom_add_cc_temp_1;
output 	rom_add_cc_temp_2;
output 	rom_add_cc_temp_3;
output 	rom_add_cc_temp_4;
output 	rom_add_cc_temp_5;
output 	rom_add_cs_6;
output 	rom_add_cs_7;
output 	rom_add_cc_temp_6;
output 	rom_add_cc_temp_7;
output 	rom_add_f_0;
output 	rom_add_f_1;
output 	rom_add_f_2;
output 	rom_add_f_3;
output 	rom_add_f_4;
output 	rom_add_f_5;
output 	rom_add_f_6;
output 	rom_add_f_7;
input 	result_a_28;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_12;
input 	pipeline_dffe_13;
input 	pipeline_dffe_14;
input 	pipeline_dffe_15;
input 	pipeline_dffe_0;
input 	pipeline_dffe_1;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;


dffeas \rom_add_cc_temp[0] (
	.clk(clk),
	.d(pipeline_dffe_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_cc_temp_0),
	.prn(vcc));
defparam \rom_add_cc_temp[0] .is_wysiwyg = "true";
defparam \rom_add_cc_temp[0] .power_up = "low";

dffeas \rom_add_cc_temp[1] (
	.clk(clk),
	.d(pipeline_dffe_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_cc_temp_1),
	.prn(vcc));
defparam \rom_add_cc_temp[1] .is_wysiwyg = "true";
defparam \rom_add_cc_temp[1] .power_up = "low";

dffeas \rom_add_cc_temp[2] (
	.clk(clk),
	.d(pipeline_dffe_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_cc_temp_2),
	.prn(vcc));
defparam \rom_add_cc_temp[2] .is_wysiwyg = "true";
defparam \rom_add_cc_temp[2] .power_up = "low";

dffeas \rom_add_cc_temp[3] (
	.clk(clk),
	.d(pipeline_dffe_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_cc_temp_3),
	.prn(vcc));
defparam \rom_add_cc_temp[3] .is_wysiwyg = "true";
defparam \rom_add_cc_temp[3] .power_up = "low";

dffeas \rom_add_cc_temp[4] (
	.clk(clk),
	.d(pipeline_dffe_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_cc_temp_4),
	.prn(vcc));
defparam \rom_add_cc_temp[4] .is_wysiwyg = "true";
defparam \rom_add_cc_temp[4] .power_up = "low";

dffeas \rom_add_cc_temp[5] (
	.clk(clk),
	.d(pipeline_dffe_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_cc_temp_5),
	.prn(vcc));
defparam \rom_add_cc_temp[5] .is_wysiwyg = "true";
defparam \rom_add_cc_temp[5] .power_up = "low";

dffeas \rom_add_cs[6] (
	.clk(clk),
	.d(pipeline_dffe_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_cs_6),
	.prn(vcc));
defparam \rom_add_cs[6] .is_wysiwyg = "true";
defparam \rom_add_cs[6] .power_up = "low";

dffeas \rom_add_cs[7] (
	.clk(clk),
	.d(pipeline_dffe_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_cs_7),
	.prn(vcc));
defparam \rom_add_cs[7] .is_wysiwyg = "true";
defparam \rom_add_cs[7] .power_up = "low";

dffeas \rom_add_cc_temp[6] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_cc_temp_6),
	.prn(vcc));
defparam \rom_add_cc_temp[6] .is_wysiwyg = "true";
defparam \rom_add_cc_temp[6] .power_up = "low";

dffeas \rom_add_cc_temp[7] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_cc_temp_7),
	.prn(vcc));
defparam \rom_add_cc_temp[7] .is_wysiwyg = "true";
defparam \rom_add_cc_temp[7] .power_up = "low";

dffeas \rom_add_f[0] (
	.clk(clk),
	.d(pipeline_dffe_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_f_0),
	.prn(vcc));
defparam \rom_add_f[0] .is_wysiwyg = "true";
defparam \rom_add_f[0] .power_up = "low";

dffeas \rom_add_f[1] (
	.clk(clk),
	.d(pipeline_dffe_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_f_1),
	.prn(vcc));
defparam \rom_add_f[1] .is_wysiwyg = "true";
defparam \rom_add_f[1] .power_up = "low";

dffeas \rom_add_f[2] (
	.clk(clk),
	.d(pipeline_dffe_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_f_2),
	.prn(vcc));
defparam \rom_add_f[2] .is_wysiwyg = "true";
defparam \rom_add_f[2] .power_up = "low";

dffeas \rom_add_f[3] (
	.clk(clk),
	.d(pipeline_dffe_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_f_3),
	.prn(vcc));
defparam \rom_add_f[3] .is_wysiwyg = "true";
defparam \rom_add_f[3] .power_up = "low";

dffeas \rom_add_f[4] (
	.clk(clk),
	.d(pipeline_dffe_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_f_4),
	.prn(vcc));
defparam \rom_add_f[4] .is_wysiwyg = "true";
defparam \rom_add_f[4] .power_up = "low";

dffeas \rom_add_f[5] (
	.clk(clk),
	.d(pipeline_dffe_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_f_5),
	.prn(vcc));
defparam \rom_add_f[5] .is_wysiwyg = "true";
defparam \rom_add_f[5] .power_up = "low";

dffeas \rom_add_f[6] (
	.clk(clk),
	.d(pipeline_dffe_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_f_6),
	.prn(vcc));
defparam \rom_add_f[6] .is_wysiwyg = "true";
defparam \rom_add_f[6] .power_up = "low";

dffeas \rom_add_f[7] (
	.clk(clk),
	.d(pipeline_dffe_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(rom_add_f_7),
	.prn(vcc));
defparam \rom_add_f[7] .is_wysiwyg = "true";
defparam \rom_add_f[7] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

endmodule

module sine_asj_nco_as_m_cen (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	q_a_10,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	q_a_16,
	q_a_17,
	q_a_18,
	q_a_19,
	q_a_20,
	q_a_21,
	q_a_22,
	q_a_23,
	rom_add_f_0,
	rom_add_f_1,
	rom_add_f_2,
	rom_add_f_3,
	rom_add_f_4,
	rom_add_f_5,
	rom_add_f_6,
	rom_add_f_7,
	clk,
	clken)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
output 	q_a_10;
output 	q_a_11;
output 	q_a_12;
output 	q_a_13;
output 	q_a_14;
output 	q_a_15;
output 	q_a_16;
output 	q_a_17;
output 	q_a_18;
output 	q_a_19;
output 	q_a_20;
output 	q_a_21;
output 	q_a_22;
output 	q_a_23;
input 	rom_add_f_0;
input 	rom_add_f_1;
input 	rom_add_f_2;
input 	rom_add_f_3;
input 	rom_add_f_4;
input 	rom_add_f_5;
input 	rom_add_f_6;
input 	rom_add_f_7;
input 	clk;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_altsyncram_1 altsyncram_component0(
	.q_a({q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.address_a({rom_add_f_7,rom_add_f_6,rom_add_f_5,rom_add_f_4,rom_add_f_3,rom_add_f_2,rom_add_f_1,rom_add_f_0}),
	.clock0(clk),
	.clocken0(clken));

endmodule

module sine_altsyncram_1 (
	q_a,
	address_a,
	clock0,
	clocken0)/* synthesis synthesis_greybox=1 */;
output 	[23:0] q_a;
input 	[7:0] address_a;
input 	clock0;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_altsyncram_m5g1 auto_generated(
	.q_a({q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0),
	.clocken0(clocken0));

endmodule

module sine_altsyncram_m5g1 (
	q_a,
	address_a,
	clock0,
	clocken0)/* synthesis synthesis_greybox=1 */;
output 	[23:0] q_a;
input 	[7:0] address_a;
input 	clock0;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 24;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "FFF000007FFE007FC01FC07F03F03F07E0F83E0F07C3E1E0F0F0787878787878";

cyclonev_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 24;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "FFFFFFFF8000007FFFE0007FFC003FF800FFC00FF803FE00FF007F807F807F80";

cyclonev_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 24;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "AAAAAAAAAAAAAAD55555552AAAAA955555AAAAA55556AAAA55552AAAD5552AAA";

cyclonev_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 24;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "33333333333333666666664CCCCCD999993333366664CCCC9999B33366664CCC";

cyclonev_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 24;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "3C3C3C3C3C3C3C7878787870F0F0E1E1E1C3C3C787870F0F1E1E3C3C787870F0";

cyclonev_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 24;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "6A956A956A956AD52AD52AD5AA55AB54AB56A952AD52A55AB54A956AD52AD5AA";

cyclonev_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 24;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "4CD9B3264CD9B3664C99B366CC993266CD9B3264C99B366CD993264C99B366CC";

cyclonev_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 24;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "70E1C3C78F1E3C7870E1C3870F1E3C78F1E3C3870E1C3870E1E3C78F1E3C78F0";

cyclonev_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "rom";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "clock0";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 24;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "D5AB56AD5AB56AD52A54A952A54A952A54A956AD5AB56AD5AB56AD5AB56AD5AA";

cyclonev_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "rom";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "clock0";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 24;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "3398CE63398CE63319CC67319CC67319CC67319CC67319CC67319CC67319CC66";

cyclonev_ram_block ram_block1a10(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "rom";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "clock0";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 24;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "5AD294B5AD294B5A5296B5A5296B5A5296B5A5296B5A5296B5A5296B5A5296B4";

cyclonev_ram_block ram_block1a11(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "rom";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "clock0";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 24;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "631CE739CE318C639CE739C6318C639CE739C6318C639CE739C6318C639CE738";

cyclonev_ram_block ram_block1a12(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "rom";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "clock0";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 24;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "7C1F07C1F03E0F83E0F83E07C1F07C1F07C1F83E0F83E0F83E07C1F07C1F07C0";

cyclonev_ram_block ram_block1a13(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "rom";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "clock0";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 24;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "801FF801FFC00FFC00FFC007FE007FE007FE003FF003FF003FF801FF801FF800";

cyclonev_ram_block ram_block1a14(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "rom";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "clock0";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 24;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "001FFFFE00000FFFFF000007FFFF800007FFFFC00003FFFFC00001FFFFE00000";

cyclonev_ram_block ram_block1a15(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "rom";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "clock0";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 24;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000";

cyclonev_ram_block ram_block1a16(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk0_output_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "rom";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "clock0";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 24;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = "FFE000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000";

cyclonev_ram_block ram_block1a17(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk0_output_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "rom";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "clock0";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 24;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a18(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk0_output_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "rom";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "clock0";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 24;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a19(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk0_output_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "rom";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "clock0";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 24;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a20(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.clk0_output_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "rom";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "clock0";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 24;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a21(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.clk0_output_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "rom";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "clock0";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 24;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a22(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.clk0_output_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "rom";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "clock0";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 24;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a23(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.clk0_output_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "sine_nco_ii_0_sin_f.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0122|altsyncram:altsyncram_component0|altsyncram_m5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "rom";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "clock0";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 24;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000";

endmodule

module sine_asj_nco_as_m_cen_1 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	q_a_10,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	q_a_16,
	q_a_17,
	q_a_18,
	q_a_19,
	q_a_20,
	q_a_21,
	q_a_22,
	q_a_23,
	rom_add_f_0,
	rom_add_f_1,
	rom_add_f_2,
	rom_add_f_3,
	rom_add_f_4,
	rom_add_f_5,
	rom_add_f_6,
	rom_add_f_7,
	clk,
	clken)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_8;
output 	q_a_9;
output 	q_a_10;
output 	q_a_11;
output 	q_a_12;
output 	q_a_13;
output 	q_a_14;
output 	q_a_15;
output 	q_a_16;
output 	q_a_17;
output 	q_a_18;
output 	q_a_19;
output 	q_a_20;
output 	q_a_21;
output 	q_a_22;
output 	q_a_23;
input 	rom_add_f_0;
input 	rom_add_f_1;
input 	rom_add_f_2;
input 	rom_add_f_3;
input 	rom_add_f_4;
input 	rom_add_f_5;
input 	rom_add_f_6;
input 	rom_add_f_7;
input 	clk;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_altsyncram_2 altsyncram_component0(
	.q_a({q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.address_a({rom_add_f_7,rom_add_f_6,rom_add_f_5,rom_add_f_4,rom_add_f_3,rom_add_f_2,rom_add_f_1,rom_add_f_0}),
	.clock0(clk),
	.clocken0(clken));

endmodule

module sine_altsyncram_2 (
	q_a,
	address_a,
	clock0,
	clocken0)/* synthesis synthesis_greybox=1 */;
output 	[23:0] q_a;
input 	[7:0] address_a;
input 	clock0;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_altsyncram_h5g1 auto_generated(
	.q_a({q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0),
	.clocken0(clocken0));

endmodule

module sine_altsyncram_h5g1 (
	q_a,
	address_a,
	clock0,
	clocken0)/* synthesis synthesis_greybox=1 */;
output 	[23:0] q_a;
input 	[7:0] address_a;
input 	clock0;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 24;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "32ACC03354CFF32ACC03256C7E34B67FE6AB701C949801B54C7C65523F8D558F";

cyclonev_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 24;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "3CC96A96CC3FFC336956931C0038DB5552670FE0E6D2AB6CC3FF8664AAA4CC7F";

cyclonev_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 24;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "95A4D98E3C00003C719B25A9556A493331E0FFFF071CCDB6955552D26663C3FF";

cyclonev_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 24;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "739C387E03FFFFC07E1C39CE664C925A5AB5555552B5A4924CCCCE31E1E03FFF";

cyclonev_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 24;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "A52952AB555555552AB56B5AD2DA4936C9933333318C638E3C3C3E0FE01FFFFF";

cyclonev_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 24;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "9364C99933333333198CE739CE39C70E3870F0F0F07C1F81FC03FE001FFFFFFF";

cyclonev_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 24;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "70E3C7870F0F0F0F0783E0F83E07C0FE07F00FF00FFC007FFC0001FFFFFFFFFF";

cyclonev_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 24;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "0FE03F80FF00FF00FF801FF801FFC001FFF0000FFFFC000003FFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "rom";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "clock0";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 24;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "001FFF8000FFFF00007FFFF800003FFFFFF000000003FFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "rom";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "clock0";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 24;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "FFFFFF80000000FFFFFFFFF800000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a10(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "rom";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "clock0";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 24;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "FFFFFF800000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a11(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "rom";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "clock0";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 24;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a12(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "rom";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "clock0";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 24;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a13(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "rom";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "clock0";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 24;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a14(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "rom";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "clock0";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 24;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a15(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "rom";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "clock0";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 24;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a16(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk0_output_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "rom";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "clock0";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 24;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a17(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk0_output_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "rom";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "clock0";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 24;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a18(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk0_output_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "rom";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "clock0";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 24;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a19(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk0_output_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "rom";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "clock0";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 24;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a20(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.clk0_output_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "rom";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "clock0";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 24;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a21(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.clk0_output_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "rom";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "clock0";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 24;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a22(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.clk0_output_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "rom";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "clock0";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 24;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a23(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.clk0_output_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "sine_nco_ii_0_cos_f.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0123|altsyncram:altsyncram_component0|altsyncram_h5g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "rom";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "clock0";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 24;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000";

endmodule

module sine_asj_nco_as_m_dp_cen (
	q_a_0,
	q_b_0,
	q_a_1,
	q_b_1,
	q_a_2,
	q_b_2,
	q_a_3,
	q_b_3,
	q_a_4,
	q_b_4,
	q_a_5,
	q_b_5,
	q_a_6,
	q_b_6,
	q_a_7,
	q_b_7,
	q_a_8,
	q_b_8,
	q_a_9,
	q_b_9,
	q_a_10,
	q_b_10,
	q_a_11,
	q_b_11,
	q_a_12,
	q_b_12,
	q_a_13,
	q_b_13,
	q_a_14,
	q_b_14,
	q_a_15,
	q_b_15,
	q_a_16,
	q_b_16,
	q_a_17,
	q_b_17,
	q_a_18,
	q_b_18,
	q_a_19,
	q_b_19,
	q_a_20,
	q_b_20,
	q_a_21,
	q_b_21,
	q_a_22,
	q_b_22,
	q_a_23,
	q_b_23,
	rom_add_cc_temp_0,
	rom_add_cc_temp_1,
	rom_add_cc_temp_2,
	rom_add_cc_temp_3,
	rom_add_cc_temp_4,
	rom_add_cc_temp_5,
	rom_add_cs_6,
	rom_add_cs_7,
	rom_add_cc_temp_6,
	rom_add_cc_temp_7,
	GND_port,
	clk,
	clken)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_b_0;
output 	q_a_1;
output 	q_b_1;
output 	q_a_2;
output 	q_b_2;
output 	q_a_3;
output 	q_b_3;
output 	q_a_4;
output 	q_b_4;
output 	q_a_5;
output 	q_b_5;
output 	q_a_6;
output 	q_b_6;
output 	q_a_7;
output 	q_b_7;
output 	q_a_8;
output 	q_b_8;
output 	q_a_9;
output 	q_b_9;
output 	q_a_10;
output 	q_b_10;
output 	q_a_11;
output 	q_b_11;
output 	q_a_12;
output 	q_b_12;
output 	q_a_13;
output 	q_b_13;
output 	q_a_14;
output 	q_b_14;
output 	q_a_15;
output 	q_b_15;
output 	q_a_16;
output 	q_b_16;
output 	q_a_17;
output 	q_b_17;
output 	q_a_18;
output 	q_b_18;
output 	q_a_19;
output 	q_b_19;
output 	q_a_20;
output 	q_b_20;
output 	q_a_21;
output 	q_b_21;
output 	q_a_22;
output 	q_b_22;
output 	q_a_23;
output 	q_b_23;
input 	rom_add_cc_temp_0;
input 	rom_add_cc_temp_1;
input 	rom_add_cc_temp_2;
input 	rom_add_cc_temp_3;
input 	rom_add_cc_temp_4;
input 	rom_add_cc_temp_5;
input 	rom_add_cs_6;
input 	rom_add_cs_7;
input 	rom_add_cc_temp_6;
input 	rom_add_cc_temp_7;
input 	GND_port;
input 	clk;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_altsyncram_3 altsyncram_component(
	.q_a({q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.q_b({q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_b({rom_add_cc_temp_7,rom_add_cc_temp_6,rom_add_cc_temp_5,rom_add_cc_temp_4,rom_add_cc_temp_3,rom_add_cc_temp_2,rom_add_cc_temp_1,rom_add_cc_temp_0}),
	.address_a({rom_add_cs_7,rom_add_cs_6,gnd,gnd,gnd,gnd,gnd,gnd}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,GND_port}),
	.clock0(clk),
	.clocken0(clken));

endmodule

module sine_altsyncram_3 (
	q_a,
	q_b,
	address_b,
	address_a,
	data_a,
	clock0,
	clocken0)/* synthesis synthesis_greybox=1 */;
output 	[23:0] q_a;
output 	[23:0] q_b;
input 	[7:0] address_b;
input 	[7:0] address_a;
input 	[23:0] data_a;
input 	clock0;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_altsyncram_0ee2 auto_generated(
	.q_a({q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.q_b({q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_b({address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.address_a({address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0]}),
	.data_b({data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0]}),
	.clock0(clock0),
	.clocken0(clocken0));

endmodule

module sine_altsyncram_0ee2 (
	q_a,
	q_b,
	address_b,
	address_a,
	data_a,
	data_b,
	clock0,
	clocken0)/* synthesis synthesis_greybox=1 */;
output 	[23:0] q_a;
output 	[23:0] q_b;
input 	[7:0] address_b;
input 	[7:0] address_a;
input 	[23:0] data_a;
input 	[23:0] data_b;
input 	clock0;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "bidir_dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 24;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 8;
defparam ram_block1a0.port_b_data_in_clock = "clock0";
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 255;
defparam ram_block1a0.port_b_logical_ram_depth = 256;
defparam ram_block1a0.port_b_logical_ram_width = 24;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.port_b_write_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "D86D2AC330946CE7CE6C521986A96C36D86D2AC330946CE7CE6C521986A96C36";

cyclonev_ram_block ram_block1a1(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "bidir_dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 24;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 8;
defparam ram_block1a1.port_b_data_in_clock = "clock0";
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 255;
defparam ram_block1a1.port_b_logical_ram_depth = 256;
defparam ram_block1a1.port_b_logical_ram_width = 24;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.port_b_write_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "40EFBE8B12A3837ABD838A91A2FBEE04988294482237EF9D73EFD88824528232";

cyclonev_ram_block ram_block1a2(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "bidir_dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 24;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 8;
defparam ram_block1a2.port_b_data_in_clock = "clock0";
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 255;
defparam ram_block1a2.port_b_logical_ram_depth = 256;
defparam ram_block1a2.port_b_logical_ram_width = 24;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.port_b_write_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "D2DA991D50FE7CA28A7CFE157132B6960A3527D66249935D7593248CD7C958A0";

cyclonev_ram_block ram_block1a3(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "bidir_dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 24;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 8;
defparam ram_block1a3.port_b_data_in_clock = "clock0";
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 255;
defparam ram_block1a3.port_b_logical_ram_depth = 256;
defparam ram_block1a3.port_b_logical_ram_width = 24;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.port_b_write_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "1BA580A4392278FEFE3C89384A034BB0C15A3F7B4BDD870101C377A5BDF8B506";

cyclonev_ram_block ram_block1a4(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "bidir_dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 24;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 8;
defparam ram_block1a4.port_b_data_in_clock = "clock0";
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 255;
defparam ram_block1a4.port_b_logical_ram_depth = 256;
defparam ram_block1a4.port_b_logical_ram_width = 24;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.port_b_write_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "ACB30B3C18FDFA06C0BF7E3079A19A6A774CB4C3630205F93F40818D865A65DC";

cyclonev_ram_block ram_block1a5(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "bidir_dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 24;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 8;
defparam ram_block1a5.port_b_data_in_clock = "clock0";
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 255;
defparam ram_block1a5.port_b_logical_ram_depth = 256;
defparam ram_block1a5.port_b_logical_ram_width = 24;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.port_b_write_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "76936ED29B72DBE44FB69DB296ED92DC896CD12DE08D241BB049620F69166D22";

cyclonev_ram_block ram_block1a6(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "bidir_dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 24;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 8;
defparam ram_block1a6.port_b_data_in_clock = "clock0";
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 255;
defparam ram_block1a6.port_b_logical_ram_depth = 256;
defparam ram_block1a6.port_b_logical_ram_width = 24;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.port_b_write_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "AFBE548CBBE978BEFA3D2FBA6254FBEA5041AB734016874105C2D0059DAB0414";

cyclonev_ram_block ram_block1a7(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "bidir_dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 24;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 8;
defparam ram_block1a7.port_b_data_in_clock = "clock0";
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 255;
defparam ram_block1a7.port_b_logical_ram_depth = 256;
defparam ram_block1a7.port_b_logical_ram_width = 24;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.port_b_write_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "8E164C89F4E8B95AB53A2E5F2264D0E271E9B3760F1746A54AC5D1E0DD9B2F1C";

cyclonev_ram_block ram_block1a8(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "bidir_dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "clock0";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 24;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 8;
defparam ram_block1a8.port_b_data_in_clock = "clock0";
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 255;
defparam ram_block1a8.port_b_logical_ram_depth = 256;
defparam ram_block1a8.port_b_logical_ram_width = 24;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.port_b_write_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "A718F783BAD2E116D10E96BB83DE31CA58E7087C452D1EE92EF169447C21CE34";

cyclonev_ram_block ram_block1a9(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "bidir_dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "clock0";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 24;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 8;
defparam ram_block1a9.port_b_data_in_clock = "clock0";
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 255;
defparam ram_block1a9.port_b_logical_ram_depth = 256;
defparam ram_block1a9.port_b_logical_ram_width = 24;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.port_b_write_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "85522184A98FDCE44E77E32A430895427AADDE7B5670231BB1881CD5BCF76ABC";

cyclonev_ram_block ram_block1a10(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "bidir_dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "clock0";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 24;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 8;
defparam ram_block1a10.port_b_data_in_clock = "clock0";
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 255;
defparam ram_block1a10.port_b_logical_ram_depth = 256;
defparam ram_block1a10.port_b_logical_ram_width = 24;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.port_b_write_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "3FF3421B1851273459C91431B0859FF8C00CBDE4E7AED8CBA636EBCE4F7A6006";

cyclonev_ram_block ram_block1a11(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "bidir_dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "clock0";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 24;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 8;
defparam ram_block1a11.port_b_data_in_clock = "clock0";
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 255;
defparam ram_block1a11.port_b_logical_ram_depth = 256;
defparam ram_block1a11.port_b_logical_ram_width = 24;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.port_b_write_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "C22A1897D29F421AB085F297D230A8863DD5E7682D60BDE54F7A0D682DCF5778";

cyclonev_ram_block ram_block1a12(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "bidir_dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "clock0";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 24;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 8;
defparam ram_block1a12.port_b_data_in_clock = "clock0";
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 255;
defparam ram_block1a12.port_b_logical_ram_depth = 256;
defparam ram_block1a12.port_b_logical_ram_width = 24;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.port_b_write_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "FEB824032FD3E73839CF97E980483AFE0147DBFCD02C18C7C63068167FB7C500";

cyclonev_ram_block ram_block1a13(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "bidir_dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "clock0";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 24;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 8;
defparam ram_block1a13.port_b_data_in_clock = "clock0";
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 255;
defparam ram_block1a13.port_b_logical_ram_depth = 256;
defparam ram_block1a13.port_b_logical_ram_width = 24;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.port_b_write_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "54C6BD0B446B69E44F2DAC45A17AC654AB3942F4BB94961BB0D253BA5E8539AA";

cyclonev_ram_block ram_block1a14(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "bidir_dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "clock0";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 24;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 8;
defparam ram_block1a14.port_b_data_in_clock = "clock0";
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 255;
defparam ram_block1a14.port_b_logical_ram_depth = 256;
defparam ram_block1a14.port_b_logical_ram_width = 24;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.port_b_write_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "98FE69F9828665E82F4CC2833F2CFE32670196067D799A17D0B33D7CC0D301CC";

cyclonev_ram_block ram_block1a15(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "bidir_dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "clock0";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 24;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 8;
defparam ram_block1a15.port_b_data_in_clock = "clock0";
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 255;
defparam ram_block1a15.port_b_logical_ram_depth = 256;
defparam ram_block1a15.port_b_logical_ram_width = 24;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.port_b_write_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "E0FE1B5201AB9CB01A73AB0095B0FE0E1F01E4ADFE54634FE58C54FF6A4F01F0";

cyclonev_ram_block ram_block1a16(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk0_output_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "bidir_dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "clock0";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 24;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 8;
defparam ram_block1a16.port_b_data_in_clock = "clock0";
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock0";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 255;
defparam ram_block1a16.port_b_logical_ram_depth = 256;
defparam ram_block1a16.port_b_logical_ram_width = 24;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.port_b_write_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = "55AB5263FF9956C006D533FF8C95AB54AA54AD9C0066A93FF92ACC00736A54AA";

cyclonev_ram_block ram_block1a17(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk0_output_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "bidir_dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "clock0";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 24;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 8;
defparam ram_block1a17.port_b_data_in_clock = "clock0";
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock0";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 255;
defparam ram_block1a17.port_b_logical_ram_depth = 256;
defparam ram_block1a17.port_b_logical_ram_width = 24;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.port_b_write_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = "339936D6AAD2670001CC96AAD6D93398CC66C929552D98FFFE3369552926CC66";

cyclonev_ram_block ram_block1a18(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk0_output_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "bidir_dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "clock0";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 24;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 8;
defparam ram_block1a18.port_b_data_in_clock = "clock0";
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock0";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 255;
defparam ram_block1a18.port_b_logical_ram_depth = 256;
defparam ram_block1a18.port_b_logical_ram_width = 24;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.port_b_write_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = "A52DA49B331C7800003C7199B24B694A5AD25B64CCE387FFFFC38E664DB496B4";

cyclonev_ram_block ram_block1a19(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk0_output_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "bidir_dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "clock0";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 24;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 8;
defparam ram_block1a19.port_b_data_in_clock = "clock0";
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock0";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 255;
defparam ram_block1a19.port_b_logical_ram_depth = 256;
defparam ram_block1a19.port_b_logical_ram_width = 24;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.port_b_write_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = "C631C71C3C1F80000003F07871C718C639CE38E3C3E07FFFFFFC0F878E38E738";

cyclonev_ram_block ram_block1a20(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.clk0_output_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "bidir_dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "clock0";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 24;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 8;
defparam ram_block1a20.port_b_data_in_clock = "clock0";
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock0";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 255;
defparam ram_block1a20.port_b_logical_ram_depth = 256;
defparam ram_block1a20.port_b_logical_ram_width = 24;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.port_b_write_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = "F83E07E03FE0000000000FF80FC0F83E07C1F81FC01FFFFFFFFFF007F03F07C0";

cyclonev_ram_block ram_block1a21(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.clk0_output_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "bidir_dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "clock0";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 24;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 8;
defparam ram_block1a21.port_b_data_in_clock = "clock0";
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock0";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 255;
defparam ram_block1a21.port_b_logical_ram_depth = 256;
defparam ram_block1a21.port_b_logical_ram_width = 24;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.port_b_write_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = "FFC007FFC000000000000007FFC007FE003FF8003FFFFFFFFFFFFFF8003FF800";

cyclonev_ram_block ram_block1a22(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.clk0_output_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "bidir_dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "clock0";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 24;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 8;
defparam ram_block1a22.port_b_data_in_clock = "clock0";
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "clock0";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 255;
defparam ram_block1a22.port_b_logical_ram_depth = 256;
defparam ram_block1a22.port_b_logical_ram_width = 24;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.port_b_write_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = "FFFFF8000000000000000000003FFFFE000007FFFFFFFFFFFFFFFFFFFFC00000";

cyclonev_ram_block ram_block1a23(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.clk0_output_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "sine_nco_ii_0_sin_c.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_dp_cen:ux0220|altsyncram:altsyncram_component|altsyncram_0ee2:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "bidir_dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "clock0";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 24;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 8;
defparam ram_block1a23.port_b_data_in_clock = "clock0";
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "clock0";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 255;
defparam ram_block1a23.port_b_logical_ram_depth = 256;
defparam ram_block1a23.port_b_logical_ram_width = 24;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.port_b_write_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000";

endmodule

module sine_asj_nco_fxx (
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	clk,
	clken,
	reset_n,
	freq_mod_i_24,
	phi_inc_i_24,
	freq_mod_i_25,
	phi_inc_i_25,
	freq_mod_i_26,
	phi_inc_i_26,
	freq_mod_i_27,
	phi_inc_i_27,
	freq_mod_i_28,
	phi_inc_i_28,
	freq_mod_i_29,
	phi_inc_i_29,
	freq_mod_i_30,
	phi_inc_i_30,
	freq_mod_i_31,
	phi_inc_i_31,
	freq_mod_i_16,
	phi_inc_i_16,
	freq_mod_i_17,
	phi_inc_i_17,
	freq_mod_i_18,
	phi_inc_i_18,
	freq_mod_i_19,
	phi_inc_i_19,
	freq_mod_i_20,
	phi_inc_i_20,
	freq_mod_i_21,
	phi_inc_i_21,
	freq_mod_i_22,
	phi_inc_i_22,
	freq_mod_i_23,
	phi_inc_i_23,
	freq_mod_i_15,
	phi_inc_i_15,
	freq_mod_i_14,
	phi_inc_i_14,
	freq_mod_i_13,
	phi_inc_i_13,
	freq_mod_i_12,
	phi_inc_i_12,
	freq_mod_i_11,
	phi_inc_i_11,
	freq_mod_i_10,
	phi_inc_i_10,
	freq_mod_i_9,
	phi_inc_i_9,
	freq_mod_i_8,
	phi_inc_i_8,
	freq_mod_i_7,
	phi_inc_i_7,
	freq_mod_i_6,
	phi_inc_i_6,
	freq_mod_i_5,
	phi_inc_i_5,
	freq_mod_i_4,
	phi_inc_i_4,
	freq_mod_i_3,
	phi_inc_i_3,
	freq_mod_i_2,
	phi_inc_i_2,
	freq_mod_i_1,
	phi_inc_i_1,
	freq_mod_i_0,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
input 	clk;
input 	clken;
input 	reset_n;
input 	freq_mod_i_24;
input 	phi_inc_i_24;
input 	freq_mod_i_25;
input 	phi_inc_i_25;
input 	freq_mod_i_26;
input 	phi_inc_i_26;
input 	freq_mod_i_27;
input 	phi_inc_i_27;
input 	freq_mod_i_28;
input 	phi_inc_i_28;
input 	freq_mod_i_29;
input 	phi_inc_i_29;
input 	freq_mod_i_30;
input 	phi_inc_i_30;
input 	freq_mod_i_31;
input 	phi_inc_i_31;
input 	freq_mod_i_16;
input 	phi_inc_i_16;
input 	freq_mod_i_17;
input 	phi_inc_i_17;
input 	freq_mod_i_18;
input 	phi_inc_i_18;
input 	freq_mod_i_19;
input 	phi_inc_i_19;
input 	freq_mod_i_20;
input 	phi_inc_i_20;
input 	freq_mod_i_21;
input 	phi_inc_i_21;
input 	freq_mod_i_22;
input 	phi_inc_i_22;
input 	freq_mod_i_23;
input 	phi_inc_i_23;
input 	freq_mod_i_15;
input 	phi_inc_i_15;
input 	freq_mod_i_14;
input 	phi_inc_i_14;
input 	freq_mod_i_13;
input 	phi_inc_i_13;
input 	freq_mod_i_12;
input 	phi_inc_i_12;
input 	freq_mod_i_11;
input 	phi_inc_i_11;
input 	freq_mod_i_10;
input 	phi_inc_i_10;
input 	freq_mod_i_9;
input 	phi_inc_i_9;
input 	freq_mod_i_8;
input 	phi_inc_i_8;
input 	freq_mod_i_7;
input 	phi_inc_i_7;
input 	freq_mod_i_6;
input 	phi_inc_i_6;
input 	freq_mod_i_5;
input 	phi_inc_i_5;
input 	freq_mod_i_4;
input 	phi_inc_i_4;
input 	freq_mod_i_3;
input 	phi_inc_i_3;
input 	freq_mod_i_2;
input 	phi_inc_i_2;
input 	freq_mod_i_1;
input 	phi_inc_i_1;
input 	freq_mod_i_0;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_lpm_add_sub_2 acc(
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.clock(clk),
	.clken(clken),
	.reset_n(reset_n),
	.freq_mod_i_24(freq_mod_i_24),
	.phi_inc_i_24(phi_inc_i_24),
	.freq_mod_i_25(freq_mod_i_25),
	.phi_inc_i_25(phi_inc_i_25),
	.freq_mod_i_26(freq_mod_i_26),
	.phi_inc_i_26(phi_inc_i_26),
	.freq_mod_i_27(freq_mod_i_27),
	.phi_inc_i_27(phi_inc_i_27),
	.freq_mod_i_28(freq_mod_i_28),
	.phi_inc_i_28(phi_inc_i_28),
	.freq_mod_i_29(freq_mod_i_29),
	.phi_inc_i_29(phi_inc_i_29),
	.freq_mod_i_30(freq_mod_i_30),
	.phi_inc_i_30(phi_inc_i_30),
	.freq_mod_i_31(freq_mod_i_31),
	.phi_inc_i_31(phi_inc_i_31),
	.freq_mod_i_16(freq_mod_i_16),
	.phi_inc_i_16(phi_inc_i_16),
	.freq_mod_i_17(freq_mod_i_17),
	.phi_inc_i_17(phi_inc_i_17),
	.freq_mod_i_18(freq_mod_i_18),
	.phi_inc_i_18(phi_inc_i_18),
	.freq_mod_i_19(freq_mod_i_19),
	.phi_inc_i_19(phi_inc_i_19),
	.freq_mod_i_20(freq_mod_i_20),
	.phi_inc_i_20(phi_inc_i_20),
	.freq_mod_i_21(freq_mod_i_21),
	.phi_inc_i_21(phi_inc_i_21),
	.freq_mod_i_22(freq_mod_i_22),
	.phi_inc_i_22(phi_inc_i_22),
	.freq_mod_i_23(freq_mod_i_23),
	.phi_inc_i_23(phi_inc_i_23),
	.freq_mod_i_15(freq_mod_i_15),
	.phi_inc_i_15(phi_inc_i_15),
	.freq_mod_i_14(freq_mod_i_14),
	.phi_inc_i_14(phi_inc_i_14),
	.freq_mod_i_13(freq_mod_i_13),
	.phi_inc_i_13(phi_inc_i_13),
	.freq_mod_i_12(freq_mod_i_12),
	.phi_inc_i_12(phi_inc_i_12),
	.freq_mod_i_11(freq_mod_i_11),
	.phi_inc_i_11(phi_inc_i_11),
	.freq_mod_i_10(freq_mod_i_10),
	.phi_inc_i_10(phi_inc_i_10),
	.freq_mod_i_9(freq_mod_i_9),
	.phi_inc_i_9(phi_inc_i_9),
	.freq_mod_i_8(freq_mod_i_8),
	.phi_inc_i_8(phi_inc_i_8),
	.freq_mod_i_7(freq_mod_i_7),
	.phi_inc_i_7(phi_inc_i_7),
	.freq_mod_i_6(freq_mod_i_6),
	.phi_inc_i_6(phi_inc_i_6),
	.freq_mod_i_5(freq_mod_i_5),
	.phi_inc_i_5(phi_inc_i_5),
	.freq_mod_i_4(freq_mod_i_4),
	.phi_inc_i_4(phi_inc_i_4),
	.freq_mod_i_3(freq_mod_i_3),
	.phi_inc_i_3(phi_inc_i_3),
	.freq_mod_i_2(freq_mod_i_2),
	.phi_inc_i_2(phi_inc_i_2),
	.freq_mod_i_1(freq_mod_i_1),
	.phi_inc_i_1(phi_inc_i_1),
	.freq_mod_i_0(freq_mod_i_0),
	.phi_inc_i_0(phi_inc_i_0));

endmodule

module sine_lpm_add_sub_2 (
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	clock,
	clken,
	reset_n,
	freq_mod_i_24,
	phi_inc_i_24,
	freq_mod_i_25,
	phi_inc_i_25,
	freq_mod_i_26,
	phi_inc_i_26,
	freq_mod_i_27,
	phi_inc_i_27,
	freq_mod_i_28,
	phi_inc_i_28,
	freq_mod_i_29,
	phi_inc_i_29,
	freq_mod_i_30,
	phi_inc_i_30,
	freq_mod_i_31,
	phi_inc_i_31,
	freq_mod_i_16,
	phi_inc_i_16,
	freq_mod_i_17,
	phi_inc_i_17,
	freq_mod_i_18,
	phi_inc_i_18,
	freq_mod_i_19,
	phi_inc_i_19,
	freq_mod_i_20,
	phi_inc_i_20,
	freq_mod_i_21,
	phi_inc_i_21,
	freq_mod_i_22,
	phi_inc_i_22,
	freq_mod_i_23,
	phi_inc_i_23,
	freq_mod_i_15,
	phi_inc_i_15,
	freq_mod_i_14,
	phi_inc_i_14,
	freq_mod_i_13,
	phi_inc_i_13,
	freq_mod_i_12,
	phi_inc_i_12,
	freq_mod_i_11,
	phi_inc_i_11,
	freq_mod_i_10,
	phi_inc_i_10,
	freq_mod_i_9,
	phi_inc_i_9,
	freq_mod_i_8,
	phi_inc_i_8,
	freq_mod_i_7,
	phi_inc_i_7,
	freq_mod_i_6,
	phi_inc_i_6,
	freq_mod_i_5,
	phi_inc_i_5,
	freq_mod_i_4,
	phi_inc_i_4,
	freq_mod_i_3,
	phi_inc_i_3,
	freq_mod_i_2,
	phi_inc_i_2,
	freq_mod_i_1,
	phi_inc_i_1,
	freq_mod_i_0,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
input 	clock;
input 	clken;
input 	reset_n;
input 	freq_mod_i_24;
input 	phi_inc_i_24;
input 	freq_mod_i_25;
input 	phi_inc_i_25;
input 	freq_mod_i_26;
input 	phi_inc_i_26;
input 	freq_mod_i_27;
input 	phi_inc_i_27;
input 	freq_mod_i_28;
input 	phi_inc_i_28;
input 	freq_mod_i_29;
input 	phi_inc_i_29;
input 	freq_mod_i_30;
input 	phi_inc_i_30;
input 	freq_mod_i_31;
input 	phi_inc_i_31;
input 	freq_mod_i_16;
input 	phi_inc_i_16;
input 	freq_mod_i_17;
input 	phi_inc_i_17;
input 	freq_mod_i_18;
input 	phi_inc_i_18;
input 	freq_mod_i_19;
input 	phi_inc_i_19;
input 	freq_mod_i_20;
input 	phi_inc_i_20;
input 	freq_mod_i_21;
input 	phi_inc_i_21;
input 	freq_mod_i_22;
input 	phi_inc_i_22;
input 	freq_mod_i_23;
input 	phi_inc_i_23;
input 	freq_mod_i_15;
input 	phi_inc_i_15;
input 	freq_mod_i_14;
input 	phi_inc_i_14;
input 	freq_mod_i_13;
input 	phi_inc_i_13;
input 	freq_mod_i_12;
input 	phi_inc_i_12;
input 	freq_mod_i_11;
input 	phi_inc_i_11;
input 	freq_mod_i_10;
input 	phi_inc_i_10;
input 	freq_mod_i_9;
input 	phi_inc_i_9;
input 	freq_mod_i_8;
input 	phi_inc_i_8;
input 	freq_mod_i_7;
input 	phi_inc_i_7;
input 	freq_mod_i_6;
input 	phi_inc_i_6;
input 	freq_mod_i_5;
input 	phi_inc_i_5;
input 	freq_mod_i_4;
input 	phi_inc_i_4;
input 	freq_mod_i_3;
input 	phi_inc_i_3;
input 	freq_mod_i_2;
input 	phi_inc_i_2;
input 	freq_mod_i_1;
input 	phi_inc_i_1;
input 	freq_mod_i_0;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_add_sub_q0h auto_generated(
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.clock(clock),
	.clken(clken),
	.reset_n(reset_n),
	.freq_mod_i_24(freq_mod_i_24),
	.phi_inc_i_24(phi_inc_i_24),
	.freq_mod_i_25(freq_mod_i_25),
	.phi_inc_i_25(phi_inc_i_25),
	.freq_mod_i_26(freq_mod_i_26),
	.phi_inc_i_26(phi_inc_i_26),
	.freq_mod_i_27(freq_mod_i_27),
	.phi_inc_i_27(phi_inc_i_27),
	.freq_mod_i_28(freq_mod_i_28),
	.phi_inc_i_28(phi_inc_i_28),
	.freq_mod_i_29(freq_mod_i_29),
	.phi_inc_i_29(phi_inc_i_29),
	.freq_mod_i_30(freq_mod_i_30),
	.phi_inc_i_30(phi_inc_i_30),
	.freq_mod_i_31(freq_mod_i_31),
	.phi_inc_i_31(phi_inc_i_31),
	.freq_mod_i_16(freq_mod_i_16),
	.phi_inc_i_16(phi_inc_i_16),
	.freq_mod_i_17(freq_mod_i_17),
	.phi_inc_i_17(phi_inc_i_17),
	.freq_mod_i_18(freq_mod_i_18),
	.phi_inc_i_18(phi_inc_i_18),
	.freq_mod_i_19(freq_mod_i_19),
	.phi_inc_i_19(phi_inc_i_19),
	.freq_mod_i_20(freq_mod_i_20),
	.phi_inc_i_20(phi_inc_i_20),
	.freq_mod_i_21(freq_mod_i_21),
	.phi_inc_i_21(phi_inc_i_21),
	.freq_mod_i_22(freq_mod_i_22),
	.phi_inc_i_22(phi_inc_i_22),
	.freq_mod_i_23(freq_mod_i_23),
	.phi_inc_i_23(phi_inc_i_23),
	.freq_mod_i_15(freq_mod_i_15),
	.phi_inc_i_15(phi_inc_i_15),
	.freq_mod_i_14(freq_mod_i_14),
	.phi_inc_i_14(phi_inc_i_14),
	.freq_mod_i_13(freq_mod_i_13),
	.phi_inc_i_13(phi_inc_i_13),
	.freq_mod_i_12(freq_mod_i_12),
	.phi_inc_i_12(phi_inc_i_12),
	.freq_mod_i_11(freq_mod_i_11),
	.phi_inc_i_11(phi_inc_i_11),
	.freq_mod_i_10(freq_mod_i_10),
	.phi_inc_i_10(phi_inc_i_10),
	.freq_mod_i_9(freq_mod_i_9),
	.phi_inc_i_9(phi_inc_i_9),
	.freq_mod_i_8(freq_mod_i_8),
	.phi_inc_i_8(phi_inc_i_8),
	.freq_mod_i_7(freq_mod_i_7),
	.phi_inc_i_7(phi_inc_i_7),
	.freq_mod_i_6(freq_mod_i_6),
	.phi_inc_i_6(phi_inc_i_6),
	.freq_mod_i_5(freq_mod_i_5),
	.phi_inc_i_5(phi_inc_i_5),
	.freq_mod_i_4(freq_mod_i_4),
	.phi_inc_i_4(phi_inc_i_4),
	.freq_mod_i_3(freq_mod_i_3),
	.phi_inc_i_3(phi_inc_i_3),
	.freq_mod_i_2(freq_mod_i_2),
	.phi_inc_i_2(phi_inc_i_2),
	.freq_mod_i_1(freq_mod_i_1),
	.phi_inc_i_1(phi_inc_i_1),
	.freq_mod_i_0(freq_mod_i_0),
	.phi_inc_i_0(phi_inc_i_0));

endmodule

module sine_add_sub_q0h (
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	clock,
	clken,
	reset_n,
	freq_mod_i_24,
	phi_inc_i_24,
	freq_mod_i_25,
	phi_inc_i_25,
	freq_mod_i_26,
	phi_inc_i_26,
	freq_mod_i_27,
	phi_inc_i_27,
	freq_mod_i_28,
	phi_inc_i_28,
	freq_mod_i_29,
	phi_inc_i_29,
	freq_mod_i_30,
	phi_inc_i_30,
	freq_mod_i_31,
	phi_inc_i_31,
	freq_mod_i_16,
	phi_inc_i_16,
	freq_mod_i_17,
	phi_inc_i_17,
	freq_mod_i_18,
	phi_inc_i_18,
	freq_mod_i_19,
	phi_inc_i_19,
	freq_mod_i_20,
	phi_inc_i_20,
	freq_mod_i_21,
	phi_inc_i_21,
	freq_mod_i_22,
	phi_inc_i_22,
	freq_mod_i_23,
	phi_inc_i_23,
	freq_mod_i_15,
	phi_inc_i_15,
	freq_mod_i_14,
	phi_inc_i_14,
	freq_mod_i_13,
	phi_inc_i_13,
	freq_mod_i_12,
	phi_inc_i_12,
	freq_mod_i_11,
	phi_inc_i_11,
	freq_mod_i_10,
	phi_inc_i_10,
	freq_mod_i_9,
	phi_inc_i_9,
	freq_mod_i_8,
	phi_inc_i_8,
	freq_mod_i_7,
	phi_inc_i_7,
	freq_mod_i_6,
	phi_inc_i_6,
	freq_mod_i_5,
	phi_inc_i_5,
	freq_mod_i_4,
	phi_inc_i_4,
	freq_mod_i_3,
	phi_inc_i_3,
	freq_mod_i_2,
	phi_inc_i_2,
	freq_mod_i_1,
	phi_inc_i_1,
	freq_mod_i_0,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
input 	clock;
input 	clken;
input 	reset_n;
input 	freq_mod_i_24;
input 	phi_inc_i_24;
input 	freq_mod_i_25;
input 	phi_inc_i_25;
input 	freq_mod_i_26;
input 	phi_inc_i_26;
input 	freq_mod_i_27;
input 	phi_inc_i_27;
input 	freq_mod_i_28;
input 	phi_inc_i_28;
input 	freq_mod_i_29;
input 	phi_inc_i_29;
input 	freq_mod_i_30;
input 	phi_inc_i_30;
input 	freq_mod_i_31;
input 	phi_inc_i_31;
input 	freq_mod_i_16;
input 	phi_inc_i_16;
input 	freq_mod_i_17;
input 	phi_inc_i_17;
input 	freq_mod_i_18;
input 	phi_inc_i_18;
input 	freq_mod_i_19;
input 	phi_inc_i_19;
input 	freq_mod_i_20;
input 	phi_inc_i_20;
input 	freq_mod_i_21;
input 	phi_inc_i_21;
input 	freq_mod_i_22;
input 	phi_inc_i_22;
input 	freq_mod_i_23;
input 	phi_inc_i_23;
input 	freq_mod_i_15;
input 	phi_inc_i_15;
input 	freq_mod_i_14;
input 	phi_inc_i_14;
input 	freq_mod_i_13;
input 	phi_inc_i_13;
input 	freq_mod_i_12;
input 	phi_inc_i_12;
input 	freq_mod_i_11;
input 	phi_inc_i_11;
input 	freq_mod_i_10;
input 	phi_inc_i_10;
input 	freq_mod_i_9;
input 	phi_inc_i_9;
input 	freq_mod_i_8;
input 	phi_inc_i_8;
input 	freq_mod_i_7;
input 	phi_inc_i_7;
input 	freq_mod_i_6;
input 	phi_inc_i_6;
input 	freq_mod_i_5;
input 	phi_inc_i_5;
input 	freq_mod_i_4;
input 	phi_inc_i_4;
input 	freq_mod_i_3;
input 	phi_inc_i_3;
input 	freq_mod_i_2;
input 	phi_inc_i_2;
input 	freq_mod_i_1;
input 	phi_inc_i_1;
input 	freq_mod_i_0;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~126 ;
wire \op_1~122 ;
wire \op_1~118 ;
wire \op_1~114 ;
wire \op_1~110 ;
wire \op_1~106 ;
wire \op_1~102 ;
wire \op_1~98 ;
wire \op_1~94 ;
wire \op_1~90 ;
wire \op_1~86 ;
wire \op_1~82 ;
wire \op_1~78 ;
wire \op_1~74 ;
wire \op_1~70 ;
wire \op_1~66 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~50 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~6 ;
wire \op_1~9_sumout ;
wire \op_1~10 ;
wire \op_1~13_sumout ;
wire \op_1~14 ;
wire \op_1~17_sumout ;
wire \op_1~18 ;
wire \op_1~21_sumout ;
wire \op_1~22 ;
wire \op_1~25_sumout ;
wire \op_1~26 ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~73_sumout ;
wire \op_1~77_sumout ;
wire \op_1~81_sumout ;
wire \op_1~85_sumout ;
wire \op_1~89_sumout ;
wire \op_1~93_sumout ;
wire \op_1~97_sumout ;
wire \op_1~101_sumout ;
wire \op_1~105_sumout ;
wire \op_1~109_sumout ;
wire \op_1~113_sumout ;
wire \op_1~117_sumout ;
wire \op_1~121_sumout ;
wire \op_1~125_sumout ;


dffeas \pipeline_dffe[24] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_24),
	.prn(vcc));
defparam \pipeline_dffe[24] .is_wysiwyg = "true";
defparam \pipeline_dffe[24] .power_up = "low";

dffeas \pipeline_dffe[25] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_25),
	.prn(vcc));
defparam \pipeline_dffe[25] .is_wysiwyg = "true";
defparam \pipeline_dffe[25] .power_up = "low";

dffeas \pipeline_dffe[26] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_26),
	.prn(vcc));
defparam \pipeline_dffe[26] .is_wysiwyg = "true";
defparam \pipeline_dffe[26] .power_up = "low";

dffeas \pipeline_dffe[27] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_27),
	.prn(vcc));
defparam \pipeline_dffe[27] .is_wysiwyg = "true";
defparam \pipeline_dffe[27] .power_up = "low";

dffeas \pipeline_dffe[28] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_28),
	.prn(vcc));
defparam \pipeline_dffe[28] .is_wysiwyg = "true";
defparam \pipeline_dffe[28] .power_up = "low";

dffeas \pipeline_dffe[29] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_29),
	.prn(vcc));
defparam \pipeline_dffe[29] .is_wysiwyg = "true";
defparam \pipeline_dffe[29] .power_up = "low";

dffeas \pipeline_dffe[30] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_30),
	.prn(vcc));
defparam \pipeline_dffe[30] .is_wysiwyg = "true";
defparam \pipeline_dffe[30] .power_up = "low";

dffeas \pipeline_dffe[31] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_31),
	.prn(vcc));
defparam \pipeline_dffe[31] .is_wysiwyg = "true";
defparam \pipeline_dffe[31] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[18] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \pipeline_dffe[18] .is_wysiwyg = "true";
defparam \pipeline_dffe[18] .power_up = "low";

dffeas \pipeline_dffe[19] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \pipeline_dffe[19] .is_wysiwyg = "true";
defparam \pipeline_dffe[19] .power_up = "low";

dffeas \pipeline_dffe[20] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_20),
	.prn(vcc));
defparam \pipeline_dffe[20] .is_wysiwyg = "true";
defparam \pipeline_dffe[20] .power_up = "low";

dffeas \pipeline_dffe[21] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_21),
	.prn(vcc));
defparam \pipeline_dffe[21] .is_wysiwyg = "true";
defparam \pipeline_dffe[21] .power_up = "low";

dffeas \pipeline_dffe[22] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_22),
	.prn(vcc));
defparam \pipeline_dffe[22] .is_wysiwyg = "true";
defparam \pipeline_dffe[22] .power_up = "low";

dffeas \pipeline_dffe[23] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_23),
	.prn(vcc));
defparam \pipeline_dffe[23] .is_wysiwyg = "true";
defparam \pipeline_dffe[23] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~73_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~77_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~81_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~85_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~89_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~93_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~97_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~101_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~105_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~109_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~113_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~117_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~121_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~125_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

cyclonev_lcell_comb \op_1~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_0),
	.datae(gnd),
	.dataf(!phi_inc_i_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~125_sumout ),
	.cout(\op_1~126 ),
	.shareout());
defparam \op_1~125 .extended_lut = "off";
defparam \op_1~125 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~125 .shared_arith = "off";

cyclonev_lcell_comb \op_1~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_1),
	.datae(gnd),
	.dataf(!phi_inc_i_1),
	.datag(gnd),
	.cin(\op_1~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~121_sumout ),
	.cout(\op_1~122 ),
	.shareout());
defparam \op_1~121 .extended_lut = "off";
defparam \op_1~121 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~121 .shared_arith = "off";

cyclonev_lcell_comb \op_1~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_2),
	.datae(gnd),
	.dataf(!phi_inc_i_2),
	.datag(gnd),
	.cin(\op_1~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~117_sumout ),
	.cout(\op_1~118 ),
	.shareout());
defparam \op_1~117 .extended_lut = "off";
defparam \op_1~117 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~117 .shared_arith = "off";

cyclonev_lcell_comb \op_1~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_3),
	.datae(gnd),
	.dataf(!phi_inc_i_3),
	.datag(gnd),
	.cin(\op_1~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~113_sumout ),
	.cout(\op_1~114 ),
	.shareout());
defparam \op_1~113 .extended_lut = "off";
defparam \op_1~113 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~113 .shared_arith = "off";

cyclonev_lcell_comb \op_1~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_4),
	.datae(gnd),
	.dataf(!phi_inc_i_4),
	.datag(gnd),
	.cin(\op_1~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~109_sumout ),
	.cout(\op_1~110 ),
	.shareout());
defparam \op_1~109 .extended_lut = "off";
defparam \op_1~109 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~109 .shared_arith = "off";

cyclonev_lcell_comb \op_1~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_5),
	.datae(gnd),
	.dataf(!phi_inc_i_5),
	.datag(gnd),
	.cin(\op_1~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~105_sumout ),
	.cout(\op_1~106 ),
	.shareout());
defparam \op_1~105 .extended_lut = "off";
defparam \op_1~105 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~105 .shared_arith = "off";

cyclonev_lcell_comb \op_1~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_6),
	.datae(gnd),
	.dataf(!phi_inc_i_6),
	.datag(gnd),
	.cin(\op_1~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~101_sumout ),
	.cout(\op_1~102 ),
	.shareout());
defparam \op_1~101 .extended_lut = "off";
defparam \op_1~101 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~101 .shared_arith = "off";

cyclonev_lcell_comb \op_1~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_7),
	.datae(gnd),
	.dataf(!phi_inc_i_7),
	.datag(gnd),
	.cin(\op_1~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~97_sumout ),
	.cout(\op_1~98 ),
	.shareout());
defparam \op_1~97 .extended_lut = "off";
defparam \op_1~97 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~97 .shared_arith = "off";

cyclonev_lcell_comb \op_1~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_8),
	.datae(gnd),
	.dataf(!phi_inc_i_8),
	.datag(gnd),
	.cin(\op_1~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~93_sumout ),
	.cout(\op_1~94 ),
	.shareout());
defparam \op_1~93 .extended_lut = "off";
defparam \op_1~93 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~93 .shared_arith = "off";

cyclonev_lcell_comb \op_1~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_9),
	.datae(gnd),
	.dataf(!phi_inc_i_9),
	.datag(gnd),
	.cin(\op_1~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~89_sumout ),
	.cout(\op_1~90 ),
	.shareout());
defparam \op_1~89 .extended_lut = "off";
defparam \op_1~89 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~89 .shared_arith = "off";

cyclonev_lcell_comb \op_1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_10),
	.datae(gnd),
	.dataf(!phi_inc_i_10),
	.datag(gnd),
	.cin(\op_1~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~85_sumout ),
	.cout(\op_1~86 ),
	.shareout());
defparam \op_1~85 .extended_lut = "off";
defparam \op_1~85 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~85 .shared_arith = "off";

cyclonev_lcell_comb \op_1~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_11),
	.datae(gnd),
	.dataf(!phi_inc_i_11),
	.datag(gnd),
	.cin(\op_1~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~81_sumout ),
	.cout(\op_1~82 ),
	.shareout());
defparam \op_1~81 .extended_lut = "off";
defparam \op_1~81 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~81 .shared_arith = "off";

cyclonev_lcell_comb \op_1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_12),
	.datae(gnd),
	.dataf(!phi_inc_i_12),
	.datag(gnd),
	.cin(\op_1~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~77_sumout ),
	.cout(\op_1~78 ),
	.shareout());
defparam \op_1~77 .extended_lut = "off";
defparam \op_1~77 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~77 .shared_arith = "off";

cyclonev_lcell_comb \op_1~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_13),
	.datae(gnd),
	.dataf(!phi_inc_i_13),
	.datag(gnd),
	.cin(\op_1~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~73_sumout ),
	.cout(\op_1~74 ),
	.shareout());
defparam \op_1~73 .extended_lut = "off";
defparam \op_1~73 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~73 .shared_arith = "off";

cyclonev_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_14),
	.datae(gnd),
	.dataf(!phi_inc_i_14),
	.datag(gnd),
	.cin(\op_1~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

cyclonev_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_15),
	.datae(gnd),
	.dataf(!phi_inc_i_15),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_16),
	.datae(gnd),
	.dataf(!phi_inc_i_16),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_17),
	.datae(gnd),
	.dataf(!phi_inc_i_17),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_18),
	.datae(gnd),
	.dataf(!phi_inc_i_18),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_19),
	.datae(gnd),
	.dataf(!phi_inc_i_19),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_20),
	.datae(gnd),
	.dataf(!phi_inc_i_20),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

cyclonev_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_21),
	.datae(gnd),
	.dataf(!phi_inc_i_21),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

cyclonev_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_22),
	.datae(gnd),
	.dataf(!phi_inc_i_22),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

cyclonev_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_23),
	.datae(gnd),
	.dataf(!phi_inc_i_23),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_24),
	.datae(gnd),
	.dataf(!phi_inc_i_24),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_25),
	.datae(gnd),
	.dataf(!phi_inc_i_25),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_26),
	.datae(gnd),
	.dataf(!phi_inc_i_26),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_27),
	.datae(gnd),
	.dataf(!phi_inc_i_27),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_28),
	.datae(gnd),
	.dataf(!phi_inc_i_28),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_29),
	.datae(gnd),
	.dataf(!phi_inc_i_29),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_30),
	.datae(gnd),
	.dataf(!phi_inc_i_30),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_31),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

endmodule

module sine_asj_nco_isdr (
	data_ready1,
	clk,
	clken,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	data_ready1;
input 	clk;
input 	clken;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lpm_counter_component|auto_generated|counter_reg_bit[3]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[2]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[1]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[0]~q ;
wire \data_ready~0_combout ;


sine_lpm_counter_1 lpm_counter_component(
	.counter_reg_bit_3(\lpm_counter_component|auto_generated|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\lpm_counter_component|auto_generated|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\lpm_counter_component|auto_generated|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\lpm_counter_component|auto_generated|counter_reg_bit[0]~q ),
	.clock(clk),
	.clken(clken),
	.sclr(reset_n));

dffeas data_ready(
	.clk(clk),
	.d(\data_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(data_ready1),
	.prn(vcc));
defparam data_ready.is_wysiwyg = "true";
defparam data_ready.power_up = "low";

cyclonev_lcell_comb \data_ready~0 (
	.dataa(!data_ready1),
	.datab(!clken),
	.datac(!\lpm_counter_component|auto_generated|counter_reg_bit[3]~q ),
	.datad(!\lpm_counter_component|auto_generated|counter_reg_bit[2]~q ),
	.datae(!\lpm_counter_component|auto_generated|counter_reg_bit[1]~q ),
	.dataf(!\lpm_counter_component|auto_generated|counter_reg_bit[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_ready~0 .extended_lut = "off";
defparam \data_ready~0 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \data_ready~0 .shared_arith = "off";

endmodule

module sine_lpm_counter_1 (
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	clock,
	clken,
	sclr)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	clock;
input 	clken;
input 	sclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_cntr_ski auto_generated(
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.clock(clock),
	.clken(clken),
	.sclr(sclr));

endmodule

module sine_cntr_ski (
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	clock,
	clken,
	sclr)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	clock;
input 	clken;
input 	sclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita0~sumout ;


dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

endmodule

module sine_asj_nco_mob_w (
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	dffe47,
	result_a_28,
	dffe24,
	dffe35,
	dffe48,
	dffe25,
	dffe26,
	dffe27,
	dffe28,
	dffe29,
	dffe30,
	dffe31,
	dffe32,
	dffe33,
	dffe34,
	dffe36,
	dffe37,
	dffe38,
	dffe39,
	dffe40,
	dffe41,
	dffe42,
	dffe43,
	dffe44,
	dffe45,
	dffe46,
	clk,
	clken,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
input 	dffe47;
input 	result_a_28;
input 	dffe24;
input 	dffe35;
input 	dffe48;
input 	dffe25;
input 	dffe26;
input 	dffe27;
input 	dffe28;
input 	dffe29;
input 	dffe30;
input 	dffe31;
input 	dffe32;
input 	dffe33;
input 	dffe34;
input 	dffe36;
input 	dffe37;
input 	dffe38;
input 	dffe39;
input 	dffe40;
input 	dffe41;
input 	dffe42;
input 	dffe43;
input 	dffe44;
input 	dffe45;
input 	dffe46;
input 	clk;
input 	clken;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_tmp[23]~q ;
wire \data_tmp[0]~q ;
wire \is_zero~q ;
wire \data_tmp[1]~q ;
wire \data_tmp[2]~q ;
wire \data_tmp[3]~q ;
wire \data_tmp[4]~q ;
wire \data_tmp[5]~q ;
wire \data_tmp[6]~q ;
wire \data_tmp[7]~q ;
wire \data_tmp[8]~q ;
wire \data_tmp[9]~q ;
wire \data_tmp[10]~q ;
wire \data_tmp[11]~q ;
wire \data_tmp[12]~q ;
wire \data_tmp[13]~q ;
wire \data_tmp[14]~q ;
wire \data_tmp[15]~q ;
wire \data_tmp[16]~q ;
wire \data_tmp[17]~q ;
wire \data_tmp[18]~q ;
wire \data_tmp[19]~q ;
wire \data_tmp[20]~q ;
wire \data_tmp[21]~q ;
wire \data_tmp[22]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \Equal0~3_combout ;
wire \Equal0~4_combout ;


sine_lpm_add_sub_3 lpm_add_sub_component(
	.data_tmp_23(\data_tmp[23]~q ),
	.data_tmp_0(\data_tmp[0]~q ),
	.is_zero(\is_zero~q ),
	.data_tmp_1(\data_tmp[1]~q ),
	.data_tmp_2(\data_tmp[2]~q ),
	.data_tmp_3(\data_tmp[3]~q ),
	.data_tmp_4(\data_tmp[4]~q ),
	.data_tmp_5(\data_tmp[5]~q ),
	.data_tmp_6(\data_tmp[6]~q ),
	.data_tmp_7(\data_tmp[7]~q ),
	.data_tmp_8(\data_tmp[8]~q ),
	.data_tmp_9(\data_tmp[9]~q ),
	.data_tmp_10(\data_tmp[10]~q ),
	.data_tmp_11(\data_tmp[11]~q ),
	.data_tmp_12(\data_tmp[12]~q ),
	.data_tmp_13(\data_tmp[13]~q ),
	.data_tmp_14(\data_tmp[14]~q ),
	.data_tmp_15(\data_tmp[15]~q ),
	.data_tmp_16(\data_tmp[16]~q ),
	.data_tmp_17(\data_tmp[17]~q ),
	.data_tmp_18(\data_tmp[18]~q ),
	.data_tmp_19(\data_tmp[19]~q ),
	.data_tmp_20(\data_tmp[20]~q ),
	.data_tmp_21(\data_tmp[21]~q ),
	.data_tmp_22(\data_tmp[22]~q ),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.clock(clk),
	.clken(clken));

dffeas \data_tmp[23] (
	.clk(clk),
	.d(dffe47),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[23]~q ),
	.prn(vcc));
defparam \data_tmp[23] .is_wysiwyg = "true";
defparam \data_tmp[23] .power_up = "low";

dffeas \data_tmp[0] (
	.clk(clk),
	.d(dffe24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[0]~q ),
	.prn(vcc));
defparam \data_tmp[0] .is_wysiwyg = "true";
defparam \data_tmp[0] .power_up = "low";

dffeas is_zero(
	.clk(clk),
	.d(\Equal0~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\is_zero~q ),
	.prn(vcc));
defparam is_zero.is_wysiwyg = "true";
defparam is_zero.power_up = "low";

dffeas \data_tmp[1] (
	.clk(clk),
	.d(dffe25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[1]~q ),
	.prn(vcc));
defparam \data_tmp[1] .is_wysiwyg = "true";
defparam \data_tmp[1] .power_up = "low";

dffeas \data_tmp[2] (
	.clk(clk),
	.d(dffe26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[2]~q ),
	.prn(vcc));
defparam \data_tmp[2] .is_wysiwyg = "true";
defparam \data_tmp[2] .power_up = "low";

dffeas \data_tmp[3] (
	.clk(clk),
	.d(dffe27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[3]~q ),
	.prn(vcc));
defparam \data_tmp[3] .is_wysiwyg = "true";
defparam \data_tmp[3] .power_up = "low";

dffeas \data_tmp[4] (
	.clk(clk),
	.d(dffe28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[4]~q ),
	.prn(vcc));
defparam \data_tmp[4] .is_wysiwyg = "true";
defparam \data_tmp[4] .power_up = "low";

dffeas \data_tmp[5] (
	.clk(clk),
	.d(dffe29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[5]~q ),
	.prn(vcc));
defparam \data_tmp[5] .is_wysiwyg = "true";
defparam \data_tmp[5] .power_up = "low";

dffeas \data_tmp[6] (
	.clk(clk),
	.d(dffe30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[6]~q ),
	.prn(vcc));
defparam \data_tmp[6] .is_wysiwyg = "true";
defparam \data_tmp[6] .power_up = "low";

dffeas \data_tmp[7] (
	.clk(clk),
	.d(dffe31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[7]~q ),
	.prn(vcc));
defparam \data_tmp[7] .is_wysiwyg = "true";
defparam \data_tmp[7] .power_up = "low";

dffeas \data_tmp[8] (
	.clk(clk),
	.d(dffe32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[8]~q ),
	.prn(vcc));
defparam \data_tmp[8] .is_wysiwyg = "true";
defparam \data_tmp[8] .power_up = "low";

dffeas \data_tmp[9] (
	.clk(clk),
	.d(dffe33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[9]~q ),
	.prn(vcc));
defparam \data_tmp[9] .is_wysiwyg = "true";
defparam \data_tmp[9] .power_up = "low";

dffeas \data_tmp[10] (
	.clk(clk),
	.d(dffe34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[10]~q ),
	.prn(vcc));
defparam \data_tmp[10] .is_wysiwyg = "true";
defparam \data_tmp[10] .power_up = "low";

dffeas \data_tmp[11] (
	.clk(clk),
	.d(dffe35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[11]~q ),
	.prn(vcc));
defparam \data_tmp[11] .is_wysiwyg = "true";
defparam \data_tmp[11] .power_up = "low";

dffeas \data_tmp[12] (
	.clk(clk),
	.d(dffe36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[12]~q ),
	.prn(vcc));
defparam \data_tmp[12] .is_wysiwyg = "true";
defparam \data_tmp[12] .power_up = "low";

dffeas \data_tmp[13] (
	.clk(clk),
	.d(dffe37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[13]~q ),
	.prn(vcc));
defparam \data_tmp[13] .is_wysiwyg = "true";
defparam \data_tmp[13] .power_up = "low";

dffeas \data_tmp[14] (
	.clk(clk),
	.d(dffe38),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[14]~q ),
	.prn(vcc));
defparam \data_tmp[14] .is_wysiwyg = "true";
defparam \data_tmp[14] .power_up = "low";

dffeas \data_tmp[15] (
	.clk(clk),
	.d(dffe39),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[15]~q ),
	.prn(vcc));
defparam \data_tmp[15] .is_wysiwyg = "true";
defparam \data_tmp[15] .power_up = "low";

dffeas \data_tmp[16] (
	.clk(clk),
	.d(dffe40),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[16]~q ),
	.prn(vcc));
defparam \data_tmp[16] .is_wysiwyg = "true";
defparam \data_tmp[16] .power_up = "low";

dffeas \data_tmp[17] (
	.clk(clk),
	.d(dffe41),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[17]~q ),
	.prn(vcc));
defparam \data_tmp[17] .is_wysiwyg = "true";
defparam \data_tmp[17] .power_up = "low";

dffeas \data_tmp[18] (
	.clk(clk),
	.d(dffe42),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[18]~q ),
	.prn(vcc));
defparam \data_tmp[18] .is_wysiwyg = "true";
defparam \data_tmp[18] .power_up = "low";

dffeas \data_tmp[19] (
	.clk(clk),
	.d(dffe43),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[19]~q ),
	.prn(vcc));
defparam \data_tmp[19] .is_wysiwyg = "true";
defparam \data_tmp[19] .power_up = "low";

dffeas \data_tmp[20] (
	.clk(clk),
	.d(dffe44),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[20]~q ),
	.prn(vcc));
defparam \data_tmp[20] .is_wysiwyg = "true";
defparam \data_tmp[20] .power_up = "low";

dffeas \data_tmp[21] (
	.clk(clk),
	.d(dffe45),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[21]~q ),
	.prn(vcc));
defparam \data_tmp[21] .is_wysiwyg = "true";
defparam \data_tmp[21] .power_up = "low";

dffeas \data_tmp[22] (
	.clk(clk),
	.d(dffe46),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\data_tmp[22]~q ),
	.prn(vcc));
defparam \data_tmp[22] .is_wysiwyg = "true";
defparam \data_tmp[22] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!dffe24),
	.datab(!dffe25),
	.datac(!dffe26),
	.datad(!dffe27),
	.datae(!dffe28),
	.dataf(!dffe29),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!dffe30),
	.datab(!dffe31),
	.datac(!dffe32),
	.datad(!dffe33),
	.datae(!dffe34),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~2 (
	.dataa(!dffe36),
	.datab(!dffe37),
	.datac(!dffe38),
	.datad(!dffe39),
	.datae(!dffe40),
	.dataf(!dffe41),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~2 .extended_lut = "off";
defparam \Equal0~2 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~3 (
	.dataa(!dffe47),
	.datab(!dffe42),
	.datac(!dffe43),
	.datad(!dffe44),
	.datae(!dffe45),
	.dataf(!dffe46),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~3 .extended_lut = "off";
defparam \Equal0~3 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal0~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~4 (
	.dataa(!dffe35),
	.datab(!dffe48),
	.datac(!\Equal0~0_combout ),
	.datad(!\Equal0~1_combout ),
	.datae(!\Equal0~2_combout ),
	.dataf(!\Equal0~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~4 .extended_lut = "off";
defparam \Equal0~4 .lut_mask = 64'hFFFFFFFFFFFFFFF7;
defparam \Equal0~4 .shared_arith = "off";

endmodule

module sine_lpm_add_sub_3 (
	data_tmp_23,
	data_tmp_0,
	is_zero,
	data_tmp_1,
	data_tmp_2,
	data_tmp_3,
	data_tmp_4,
	data_tmp_5,
	data_tmp_6,
	data_tmp_7,
	data_tmp_8,
	data_tmp_9,
	data_tmp_10,
	data_tmp_11,
	data_tmp_12,
	data_tmp_13,
	data_tmp_14,
	data_tmp_15,
	data_tmp_16,
	data_tmp_17,
	data_tmp_18,
	data_tmp_19,
	data_tmp_20,
	data_tmp_21,
	data_tmp_22,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	clock,
	clken)/* synthesis synthesis_greybox=1 */;
input 	data_tmp_23;
input 	data_tmp_0;
input 	is_zero;
input 	data_tmp_1;
input 	data_tmp_2;
input 	data_tmp_3;
input 	data_tmp_4;
input 	data_tmp_5;
input 	data_tmp_6;
input 	data_tmp_7;
input 	data_tmp_8;
input 	data_tmp_9;
input 	data_tmp_10;
input 	data_tmp_11;
input 	data_tmp_12;
input 	data_tmp_13;
input 	data_tmp_14;
input 	data_tmp_15;
input 	data_tmp_16;
input 	data_tmp_17;
input 	data_tmp_18;
input 	data_tmp_19;
input 	data_tmp_20;
input 	data_tmp_21;
input 	data_tmp_22;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
input 	clock;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_add_sub_4ik auto_generated(
	.data_tmp_23(data_tmp_23),
	.data_tmp_0(data_tmp_0),
	.is_zero(is_zero),
	.data_tmp_1(data_tmp_1),
	.data_tmp_2(data_tmp_2),
	.data_tmp_3(data_tmp_3),
	.data_tmp_4(data_tmp_4),
	.data_tmp_5(data_tmp_5),
	.data_tmp_6(data_tmp_6),
	.data_tmp_7(data_tmp_7),
	.data_tmp_8(data_tmp_8),
	.data_tmp_9(data_tmp_9),
	.data_tmp_10(data_tmp_10),
	.data_tmp_11(data_tmp_11),
	.data_tmp_12(data_tmp_12),
	.data_tmp_13(data_tmp_13),
	.data_tmp_14(data_tmp_14),
	.data_tmp_15(data_tmp_15),
	.data_tmp_16(data_tmp_16),
	.data_tmp_17(data_tmp_17),
	.data_tmp_18(data_tmp_18),
	.data_tmp_19(data_tmp_19),
	.data_tmp_20(data_tmp_20),
	.data_tmp_21(data_tmp_21),
	.data_tmp_22(data_tmp_22),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.clock(clock),
	.clken(clken));

endmodule

module sine_add_sub_4ik (
	data_tmp_23,
	data_tmp_0,
	is_zero,
	data_tmp_1,
	data_tmp_2,
	data_tmp_3,
	data_tmp_4,
	data_tmp_5,
	data_tmp_6,
	data_tmp_7,
	data_tmp_8,
	data_tmp_9,
	data_tmp_10,
	data_tmp_11,
	data_tmp_12,
	data_tmp_13,
	data_tmp_14,
	data_tmp_15,
	data_tmp_16,
	data_tmp_17,
	data_tmp_18,
	data_tmp_19,
	data_tmp_20,
	data_tmp_21,
	data_tmp_22,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	clock,
	clken)/* synthesis synthesis_greybox=1 */;
input 	data_tmp_23;
input 	data_tmp_0;
input 	is_zero;
input 	data_tmp_1;
input 	data_tmp_2;
input 	data_tmp_3;
input 	data_tmp_4;
input 	data_tmp_5;
input 	data_tmp_6;
input 	data_tmp_7;
input 	data_tmp_8;
input 	data_tmp_9;
input 	data_tmp_10;
input 	data_tmp_11;
input 	data_tmp_12;
input 	data_tmp_13;
input 	data_tmp_14;
input 	data_tmp_15;
input 	data_tmp_16;
input 	data_tmp_17;
input 	data_tmp_18;
input 	data_tmp_19;
input 	data_tmp_20;
input 	data_tmp_21;
input 	data_tmp_22;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
input 	clock;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~6 ;
wire \op_1~9_sumout ;
wire \op_1~10 ;
wire \op_1~13_sumout ;
wire \op_1~14 ;
wire \op_1~17_sumout ;
wire \op_1~18 ;
wire \op_1~21_sumout ;
wire \op_1~22 ;
wire \op_1~25_sumout ;
wire \op_1~26 ;
wire \op_1~29_sumout ;
wire \op_1~30 ;
wire \op_1~33_sumout ;
wire \op_1~34 ;
wire \op_1~37_sumout ;
wire \op_1~38 ;
wire \op_1~41_sumout ;
wire \op_1~42 ;
wire \op_1~45_sumout ;
wire \op_1~46 ;
wire \op_1~49_sumout ;
wire \op_1~50 ;
wire \op_1~53_sumout ;
wire \op_1~54 ;
wire \op_1~57_sumout ;
wire \op_1~58 ;
wire \op_1~61_sumout ;
wire \op_1~62 ;
wire \op_1~65_sumout ;
wire \op_1~66 ;
wire \op_1~69_sumout ;
wire \op_1~70 ;
wire \op_1~73_sumout ;
wire \op_1~74 ;
wire \op_1~77_sumout ;
wire \op_1~78 ;
wire \op_1~81_sumout ;
wire \op_1~82 ;
wire \op_1~85_sumout ;
wire \op_1~86 ;
wire \op_1~89_sumout ;
wire \op_1~90 ;
wire \op_1~93_sumout ;


dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[18] (
	.clk(clock),
	.d(\op_1~73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \pipeline_dffe[18] .is_wysiwyg = "true";
defparam \pipeline_dffe[18] .power_up = "low";

dffeas \pipeline_dffe[19] (
	.clk(clock),
	.d(\op_1~77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \pipeline_dffe[19] .is_wysiwyg = "true";
defparam \pipeline_dffe[19] .power_up = "low";

dffeas \pipeline_dffe[20] (
	.clk(clock),
	.d(\op_1~81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_20),
	.prn(vcc));
defparam \pipeline_dffe[20] .is_wysiwyg = "true";
defparam \pipeline_dffe[20] .power_up = "low";

dffeas \pipeline_dffe[21] (
	.clk(clock),
	.d(\op_1~85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_21),
	.prn(vcc));
defparam \pipeline_dffe[21] .is_wysiwyg = "true";
defparam \pipeline_dffe[21] .power_up = "low";

dffeas \pipeline_dffe[22] (
	.clk(clock),
	.d(\op_1~89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_22),
	.prn(vcc));
defparam \pipeline_dffe[22] .is_wysiwyg = "true";
defparam \pipeline_dffe[22] .power_up = "low";

dffeas \pipeline_dffe[23] (
	.clk(clock),
	.d(\op_1~93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_23),
	.prn(vcc));
defparam \pipeline_dffe[23] .is_wysiwyg = "true";
defparam \pipeline_dffe[23] .power_up = "low";

cyclonev_lcell_comb \op_1~1 (
	.dataa(!data_tmp_23),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_0),
	.datae(gnd),
	.dataf(!is_zero),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF55000000FF;
defparam \op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h00000000000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h00000000000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h00000000000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h00000000000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h00000000000000FF;
defparam \op_1~49 .shared_arith = "off";

cyclonev_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h00000000000000FF;
defparam \op_1~53 .shared_arith = "off";

cyclonev_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h00000000000000FF;
defparam \op_1~57 .shared_arith = "off";

cyclonev_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h00000000000000FF;
defparam \op_1~61 .shared_arith = "off";

cyclonev_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h00000000000000FF;
defparam \op_1~65 .shared_arith = "off";

cyclonev_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h00000000000000FF;
defparam \op_1~69 .shared_arith = "off";

cyclonev_lcell_comb \op_1~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~73_sumout ),
	.cout(\op_1~74 ),
	.shareout());
defparam \op_1~73 .extended_lut = "off";
defparam \op_1~73 .lut_mask = 64'h00000000000000FF;
defparam \op_1~73 .shared_arith = "off";

cyclonev_lcell_comb \op_1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_19),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~77_sumout ),
	.cout(\op_1~78 ),
	.shareout());
defparam \op_1~77 .extended_lut = "off";
defparam \op_1~77 .lut_mask = 64'h00000000000000FF;
defparam \op_1~77 .shared_arith = "off";

cyclonev_lcell_comb \op_1~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~81_sumout ),
	.cout(\op_1~82 ),
	.shareout());
defparam \op_1~81 .extended_lut = "off";
defparam \op_1~81 .lut_mask = 64'h00000000000000FF;
defparam \op_1~81 .shared_arith = "off";

cyclonev_lcell_comb \op_1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~85_sumout ),
	.cout(\op_1~86 ),
	.shareout());
defparam \op_1~85 .extended_lut = "off";
defparam \op_1~85 .lut_mask = 64'h00000000000000FF;
defparam \op_1~85 .shared_arith = "off";

cyclonev_lcell_comb \op_1~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~89_sumout ),
	.cout(\op_1~90 ),
	.shareout());
defparam \op_1~89 .extended_lut = "off";
defparam \op_1~89 .lut_mask = 64'h00000000000000FF;
defparam \op_1~89 .shared_arith = "off";

cyclonev_lcell_comb \op_1~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!data_tmp_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~93_sumout ),
	.cout(),
	.shareout());
defparam \op_1~93 .extended_lut = "off";
defparam \op_1~93 .lut_mask = 64'h00000000000000FF;
defparam \op_1~93 .shared_arith = "off";

endmodule

module sine_asj_nco_pxx (
	dxxpdo_13,
	dxxpdo_14,
	dxxpdo_15,
	dxxpdo_16,
	dxxpdo_17,
	dxxpdo_18,
	dxxpdo_19,
	dxxpdo_20,
	dxxpdo_5,
	dxxpdo_6,
	dxxpdo_7,
	dxxpdo_8,
	dxxpdo_9,
	dxxpdo_10,
	dxxpdo_11,
	dxxpdo_12,
	result_a_28,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	clk,
	clken,
	reset_n,
	phase_mod_i_8,
	phase_mod_i_9,
	phase_mod_i_10,
	phase_mod_i_11,
	phase_mod_i_12,
	phase_mod_i_13,
	phase_mod_i_14,
	phase_mod_i_15,
	phase_mod_i_0,
	phase_mod_i_1,
	phase_mod_i_2,
	phase_mod_i_3,
	phase_mod_i_4,
	phase_mod_i_5,
	phase_mod_i_6,
	phase_mod_i_7)/* synthesis synthesis_greybox=1 */;
input 	dxxpdo_13;
input 	dxxpdo_14;
input 	dxxpdo_15;
input 	dxxpdo_16;
input 	dxxpdo_17;
input 	dxxpdo_18;
input 	dxxpdo_19;
input 	dxxpdo_20;
input 	dxxpdo_5;
input 	dxxpdo_6;
input 	dxxpdo_7;
input 	dxxpdo_8;
input 	dxxpdo_9;
input 	dxxpdo_10;
input 	dxxpdo_11;
input 	dxxpdo_12;
input 	result_a_28;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
input 	clk;
input 	clken;
input 	reset_n;
input 	phase_mod_i_8;
input 	phase_mod_i_9;
input 	phase_mod_i_10;
input 	phase_mod_i_11;
input 	phase_mod_i_12;
input 	phase_mod_i_13;
input 	phase_mod_i_14;
input 	phase_mod_i_15;
input 	phase_mod_i_0;
input 	phase_mod_i_1;
input 	phase_mod_i_2;
input 	phase_mod_i_3;
input 	phase_mod_i_4;
input 	phase_mod_i_5;
input 	phase_mod_i_6;
input 	phase_mod_i_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \phi_mod_int_reg[3][8]~q ;
wire \phi_mod_int_reg[3][9]~q ;
wire \phi_mod_int_reg[3][10]~q ;
wire \phi_mod_int_reg[3][11]~q ;
wire \phi_mod_int_reg[3][12]~q ;
wire \phi_mod_int_reg[3][13]~q ;
wire \phi_mod_int_reg[3][14]~q ;
wire \phi_mod_int_reg[3][15]~q ;
wire \phi_mod_int_reg[3][0]~q ;
wire \phi_mod_int_reg[3][1]~q ;
wire \phi_mod_int_reg[3][2]~q ;
wire \phi_mod_int_reg[3][3]~q ;
wire \phi_mod_int_reg[3][4]~q ;
wire \phi_mod_int_reg[3][5]~q ;
wire \phi_mod_int_reg[3][6]~q ;
wire \phi_mod_int_reg[3][7]~q ;
wire \phi_mod_int_reg[2][8]~q ;
wire \phi_mod_int_reg[2][9]~q ;
wire \phi_mod_int_reg[2][10]~q ;
wire \phi_mod_int_reg[2][11]~q ;
wire \phi_mod_int_reg[2][12]~q ;
wire \phi_mod_int_reg[2][13]~q ;
wire \phi_mod_int_reg[2][14]~q ;
wire \phi_mod_int_reg[2][15]~q ;
wire \phi_mod_int_reg[2][0]~q ;
wire \phi_mod_int_reg[2][1]~q ;
wire \phi_mod_int_reg[2][2]~q ;
wire \phi_mod_int_reg[2][3]~q ;
wire \phi_mod_int_reg[2][4]~q ;
wire \phi_mod_int_reg[2][5]~q ;
wire \phi_mod_int_reg[2][6]~q ;
wire \phi_mod_int_reg[2][7]~q ;
wire \phi_mod_int_reg[1][8]~q ;
wire \phi_mod_int_reg[1][9]~q ;
wire \phi_mod_int_reg[1][10]~q ;
wire \phi_mod_int_reg[1][11]~q ;
wire \phi_mod_int_reg[1][12]~q ;
wire \phi_mod_int_reg[1][13]~q ;
wire \phi_mod_int_reg[1][14]~q ;
wire \phi_mod_int_reg[1][15]~q ;
wire \phi_mod_int_reg[1][0]~q ;
wire \phi_mod_int_reg[1][1]~q ;
wire \phi_mod_int_reg[1][2]~q ;
wire \phi_mod_int_reg[1][3]~q ;
wire \phi_mod_int_reg[1][4]~q ;
wire \phi_mod_int_reg[1][5]~q ;
wire \phi_mod_int_reg[1][6]~q ;
wire \phi_mod_int_reg[1][7]~q ;
wire \phi_mod_int_reg[0][8]~q ;
wire \phi_mod_int_reg[0][9]~q ;
wire \phi_mod_int_reg[0][10]~q ;
wire \phi_mod_int_reg[0][11]~q ;
wire \phi_mod_int_reg[0][12]~q ;
wire \phi_mod_int_reg[0][13]~q ;
wire \phi_mod_int_reg[0][14]~q ;
wire \phi_mod_int_reg[0][15]~q ;
wire \phi_mod_int_reg[0][0]~q ;
wire \phi_mod_int_reg[0][1]~q ;
wire \phi_mod_int_reg[0][2]~q ;
wire \phi_mod_int_reg[0][3]~q ;
wire \phi_mod_int_reg[0][4]~q ;
wire \phi_mod_int_reg[0][5]~q ;
wire \phi_mod_int_reg[0][6]~q ;
wire \phi_mod_int_reg[0][7]~q ;


sine_lpm_add_sub_4 acc(
	.dxxpdo_13(dxxpdo_13),
	.phi_mod_int_reg_8_3(\phi_mod_int_reg[3][8]~q ),
	.dxxpdo_14(dxxpdo_14),
	.phi_mod_int_reg_9_3(\phi_mod_int_reg[3][9]~q ),
	.dxxpdo_15(dxxpdo_15),
	.phi_mod_int_reg_10_3(\phi_mod_int_reg[3][10]~q ),
	.dxxpdo_16(dxxpdo_16),
	.phi_mod_int_reg_11_3(\phi_mod_int_reg[3][11]~q ),
	.dxxpdo_17(dxxpdo_17),
	.phi_mod_int_reg_12_3(\phi_mod_int_reg[3][12]~q ),
	.dxxpdo_18(dxxpdo_18),
	.phi_mod_int_reg_13_3(\phi_mod_int_reg[3][13]~q ),
	.dxxpdo_19(dxxpdo_19),
	.phi_mod_int_reg_14_3(\phi_mod_int_reg[3][14]~q ),
	.dxxpdo_20(dxxpdo_20),
	.phi_mod_int_reg_15_3(\phi_mod_int_reg[3][15]~q ),
	.dxxpdo_5(dxxpdo_5),
	.phi_mod_int_reg_0_3(\phi_mod_int_reg[3][0]~q ),
	.dxxpdo_6(dxxpdo_6),
	.phi_mod_int_reg_1_3(\phi_mod_int_reg[3][1]~q ),
	.dxxpdo_7(dxxpdo_7),
	.phi_mod_int_reg_2_3(\phi_mod_int_reg[3][2]~q ),
	.dxxpdo_8(dxxpdo_8),
	.phi_mod_int_reg_3_3(\phi_mod_int_reg[3][3]~q ),
	.dxxpdo_9(dxxpdo_9),
	.phi_mod_int_reg_4_3(\phi_mod_int_reg[3][4]~q ),
	.dxxpdo_10(dxxpdo_10),
	.phi_mod_int_reg_5_3(\phi_mod_int_reg[3][5]~q ),
	.dxxpdo_11(dxxpdo_11),
	.phi_mod_int_reg_6_3(\phi_mod_int_reg[3][6]~q ),
	.dxxpdo_12(dxxpdo_12),
	.phi_mod_int_reg_7_3(\phi_mod_int_reg[3][7]~q ),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.clock(clk),
	.clken(clken),
	.reset_n(reset_n));

dffeas \phi_mod_int_reg[3][8] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][8]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][8] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][8] .power_up = "low";

dffeas \phi_mod_int_reg[3][9] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][9]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][9] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][9] .power_up = "low";

dffeas \phi_mod_int_reg[3][10] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][10]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][10] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][10] .power_up = "low";

dffeas \phi_mod_int_reg[3][11] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][11]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][11] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][11] .power_up = "low";

dffeas \phi_mod_int_reg[3][12] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][12]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][12] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][12] .power_up = "low";

dffeas \phi_mod_int_reg[3][13] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][13]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][13] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][13] .power_up = "low";

dffeas \phi_mod_int_reg[3][14] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][14]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][14] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][14] .power_up = "low";

dffeas \phi_mod_int_reg[3][15] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][15]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][15] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][15] .power_up = "low";

dffeas \phi_mod_int_reg[3][0] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][0]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][0] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][0] .power_up = "low";

dffeas \phi_mod_int_reg[3][1] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][1]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][1] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][1] .power_up = "low";

dffeas \phi_mod_int_reg[3][2] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][2]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][2] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][2] .power_up = "low";

dffeas \phi_mod_int_reg[3][3] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][3]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][3] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][3] .power_up = "low";

dffeas \phi_mod_int_reg[3][4] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][4]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][4] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][4] .power_up = "low";

dffeas \phi_mod_int_reg[3][5] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][5]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][5] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][5] .power_up = "low";

dffeas \phi_mod_int_reg[3][6] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][6]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][6] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][6] .power_up = "low";

dffeas \phi_mod_int_reg[3][7] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[3][7]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][7] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][7] .power_up = "low";

dffeas \phi_mod_int_reg[2][8] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][8]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][8] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][8] .power_up = "low";

dffeas \phi_mod_int_reg[2][9] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][9]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][9] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][9] .power_up = "low";

dffeas \phi_mod_int_reg[2][10] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][10]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][10] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][10] .power_up = "low";

dffeas \phi_mod_int_reg[2][11] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][11]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][11] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][11] .power_up = "low";

dffeas \phi_mod_int_reg[2][12] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][12]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][12] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][12] .power_up = "low";

dffeas \phi_mod_int_reg[2][13] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][13]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][13] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][13] .power_up = "low";

dffeas \phi_mod_int_reg[2][14] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][14]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][14] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][14] .power_up = "low";

dffeas \phi_mod_int_reg[2][15] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][15]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][15] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][15] .power_up = "low";

dffeas \phi_mod_int_reg[2][0] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][0]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][0] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][0] .power_up = "low";

dffeas \phi_mod_int_reg[2][1] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][1]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][1] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][1] .power_up = "low";

dffeas \phi_mod_int_reg[2][2] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][2]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][2] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][2] .power_up = "low";

dffeas \phi_mod_int_reg[2][3] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][3]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][3] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][3] .power_up = "low";

dffeas \phi_mod_int_reg[2][4] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][4]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][4] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][4] .power_up = "low";

dffeas \phi_mod_int_reg[2][5] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][5]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][5] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][5] .power_up = "low";

dffeas \phi_mod_int_reg[2][6] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][6]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][6] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][6] .power_up = "low";

dffeas \phi_mod_int_reg[2][7] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[2][7]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][7] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][7] .power_up = "low";

dffeas \phi_mod_int_reg[1][8] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][8]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][8] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][8] .power_up = "low";

dffeas \phi_mod_int_reg[1][9] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][9]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][9] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][9] .power_up = "low";

dffeas \phi_mod_int_reg[1][10] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][10]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][10] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][10] .power_up = "low";

dffeas \phi_mod_int_reg[1][11] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][11]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][11] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][11] .power_up = "low";

dffeas \phi_mod_int_reg[1][12] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][12]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][12] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][12] .power_up = "low";

dffeas \phi_mod_int_reg[1][13] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][13]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][13] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][13] .power_up = "low";

dffeas \phi_mod_int_reg[1][14] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][14]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][14] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][14] .power_up = "low";

dffeas \phi_mod_int_reg[1][15] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][15]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][15] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][15] .power_up = "low";

dffeas \phi_mod_int_reg[1][0] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][0]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][0] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][0] .power_up = "low";

dffeas \phi_mod_int_reg[1][1] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][1]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][1] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][1] .power_up = "low";

dffeas \phi_mod_int_reg[1][2] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][2]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][2] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][2] .power_up = "low";

dffeas \phi_mod_int_reg[1][3] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][3]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][3] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][3] .power_up = "low";

dffeas \phi_mod_int_reg[1][4] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][4]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][4] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][4] .power_up = "low";

dffeas \phi_mod_int_reg[1][5] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][5]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][5] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][5] .power_up = "low";

dffeas \phi_mod_int_reg[1][6] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][6]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][6] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][6] .power_up = "low";

dffeas \phi_mod_int_reg[1][7] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[1][7]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][7] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][7] .power_up = "low";

dffeas \phi_mod_int_reg[0][8] (
	.clk(clk),
	.d(phase_mod_i_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][8]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][8] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][8] .power_up = "low";

dffeas \phi_mod_int_reg[0][9] (
	.clk(clk),
	.d(phase_mod_i_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][9]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][9] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][9] .power_up = "low";

dffeas \phi_mod_int_reg[0][10] (
	.clk(clk),
	.d(phase_mod_i_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][10]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][10] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][10] .power_up = "low";

dffeas \phi_mod_int_reg[0][11] (
	.clk(clk),
	.d(phase_mod_i_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][11]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][11] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][11] .power_up = "low";

dffeas \phi_mod_int_reg[0][12] (
	.clk(clk),
	.d(phase_mod_i_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][12]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][12] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][12] .power_up = "low";

dffeas \phi_mod_int_reg[0][13] (
	.clk(clk),
	.d(phase_mod_i_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][13]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][13] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][13] .power_up = "low";

dffeas \phi_mod_int_reg[0][14] (
	.clk(clk),
	.d(phase_mod_i_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][14]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][14] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][14] .power_up = "low";

dffeas \phi_mod_int_reg[0][15] (
	.clk(clk),
	.d(phase_mod_i_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][15]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][15] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][15] .power_up = "low";

dffeas \phi_mod_int_reg[0][0] (
	.clk(clk),
	.d(phase_mod_i_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][0]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][0] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][0] .power_up = "low";

dffeas \phi_mod_int_reg[0][1] (
	.clk(clk),
	.d(phase_mod_i_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][1]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][1] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][1] .power_up = "low";

dffeas \phi_mod_int_reg[0][2] (
	.clk(clk),
	.d(phase_mod_i_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][2]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][2] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][2] .power_up = "low";

dffeas \phi_mod_int_reg[0][3] (
	.clk(clk),
	.d(phase_mod_i_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][3]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][3] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][3] .power_up = "low";

dffeas \phi_mod_int_reg[0][4] (
	.clk(clk),
	.d(phase_mod_i_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][4]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][4] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][4] .power_up = "low";

dffeas \phi_mod_int_reg[0][5] (
	.clk(clk),
	.d(phase_mod_i_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][5]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][5] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][5] .power_up = "low";

dffeas \phi_mod_int_reg[0][6] (
	.clk(clk),
	.d(phase_mod_i_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][6]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][6] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][6] .power_up = "low";

dffeas \phi_mod_int_reg[0][7] (
	.clk(clk),
	.d(phase_mod_i_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\phi_mod_int_reg[0][7]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][7] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][7] .power_up = "low";

endmodule

module sine_lpm_add_sub_4 (
	dxxpdo_13,
	phi_mod_int_reg_8_3,
	dxxpdo_14,
	phi_mod_int_reg_9_3,
	dxxpdo_15,
	phi_mod_int_reg_10_3,
	dxxpdo_16,
	phi_mod_int_reg_11_3,
	dxxpdo_17,
	phi_mod_int_reg_12_3,
	dxxpdo_18,
	phi_mod_int_reg_13_3,
	dxxpdo_19,
	phi_mod_int_reg_14_3,
	dxxpdo_20,
	phi_mod_int_reg_15_3,
	dxxpdo_5,
	phi_mod_int_reg_0_3,
	dxxpdo_6,
	phi_mod_int_reg_1_3,
	dxxpdo_7,
	phi_mod_int_reg_2_3,
	dxxpdo_8,
	phi_mod_int_reg_3_3,
	dxxpdo_9,
	phi_mod_int_reg_4_3,
	dxxpdo_10,
	phi_mod_int_reg_5_3,
	dxxpdo_11,
	phi_mod_int_reg_6_3,
	dxxpdo_12,
	phi_mod_int_reg_7_3,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	clock,
	clken,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	dxxpdo_13;
input 	phi_mod_int_reg_8_3;
input 	dxxpdo_14;
input 	phi_mod_int_reg_9_3;
input 	dxxpdo_15;
input 	phi_mod_int_reg_10_3;
input 	dxxpdo_16;
input 	phi_mod_int_reg_11_3;
input 	dxxpdo_17;
input 	phi_mod_int_reg_12_3;
input 	dxxpdo_18;
input 	phi_mod_int_reg_13_3;
input 	dxxpdo_19;
input 	phi_mod_int_reg_14_3;
input 	dxxpdo_20;
input 	phi_mod_int_reg_15_3;
input 	dxxpdo_5;
input 	phi_mod_int_reg_0_3;
input 	dxxpdo_6;
input 	phi_mod_int_reg_1_3;
input 	dxxpdo_7;
input 	phi_mod_int_reg_2_3;
input 	dxxpdo_8;
input 	phi_mod_int_reg_3_3;
input 	dxxpdo_9;
input 	phi_mod_int_reg_4_3;
input 	dxxpdo_10;
input 	phi_mod_int_reg_5_3;
input 	dxxpdo_11;
input 	phi_mod_int_reg_6_3;
input 	dxxpdo_12;
input 	phi_mod_int_reg_7_3;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
input 	clock;
input 	clken;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_add_sub_s0h auto_generated(
	.dxxpdo_13(dxxpdo_13),
	.phi_mod_int_reg_8_3(phi_mod_int_reg_8_3),
	.dxxpdo_14(dxxpdo_14),
	.phi_mod_int_reg_9_3(phi_mod_int_reg_9_3),
	.dxxpdo_15(dxxpdo_15),
	.phi_mod_int_reg_10_3(phi_mod_int_reg_10_3),
	.dxxpdo_16(dxxpdo_16),
	.phi_mod_int_reg_11_3(phi_mod_int_reg_11_3),
	.dxxpdo_17(dxxpdo_17),
	.phi_mod_int_reg_12_3(phi_mod_int_reg_12_3),
	.dxxpdo_18(dxxpdo_18),
	.phi_mod_int_reg_13_3(phi_mod_int_reg_13_3),
	.dxxpdo_19(dxxpdo_19),
	.phi_mod_int_reg_14_3(phi_mod_int_reg_14_3),
	.dxxpdo_20(dxxpdo_20),
	.phi_mod_int_reg_15_3(phi_mod_int_reg_15_3),
	.dxxpdo_5(dxxpdo_5),
	.phi_mod_int_reg_0_3(phi_mod_int_reg_0_3),
	.dxxpdo_6(dxxpdo_6),
	.phi_mod_int_reg_1_3(phi_mod_int_reg_1_3),
	.dxxpdo_7(dxxpdo_7),
	.phi_mod_int_reg_2_3(phi_mod_int_reg_2_3),
	.dxxpdo_8(dxxpdo_8),
	.phi_mod_int_reg_3_3(phi_mod_int_reg_3_3),
	.dxxpdo_9(dxxpdo_9),
	.phi_mod_int_reg_4_3(phi_mod_int_reg_4_3),
	.dxxpdo_10(dxxpdo_10),
	.phi_mod_int_reg_5_3(phi_mod_int_reg_5_3),
	.dxxpdo_11(dxxpdo_11),
	.phi_mod_int_reg_6_3(phi_mod_int_reg_6_3),
	.dxxpdo_12(dxxpdo_12),
	.phi_mod_int_reg_7_3(phi_mod_int_reg_7_3),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.clock(clock),
	.clken(clken),
	.reset_n(reset_n));

endmodule

module sine_add_sub_s0h (
	dxxpdo_13,
	phi_mod_int_reg_8_3,
	dxxpdo_14,
	phi_mod_int_reg_9_3,
	dxxpdo_15,
	phi_mod_int_reg_10_3,
	dxxpdo_16,
	phi_mod_int_reg_11_3,
	dxxpdo_17,
	phi_mod_int_reg_12_3,
	dxxpdo_18,
	phi_mod_int_reg_13_3,
	dxxpdo_19,
	phi_mod_int_reg_14_3,
	dxxpdo_20,
	phi_mod_int_reg_15_3,
	dxxpdo_5,
	phi_mod_int_reg_0_3,
	dxxpdo_6,
	phi_mod_int_reg_1_3,
	dxxpdo_7,
	phi_mod_int_reg_2_3,
	dxxpdo_8,
	phi_mod_int_reg_3_3,
	dxxpdo_9,
	phi_mod_int_reg_4_3,
	dxxpdo_10,
	phi_mod_int_reg_5_3,
	dxxpdo_11,
	phi_mod_int_reg_6_3,
	dxxpdo_12,
	phi_mod_int_reg_7_3,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	clock,
	clken,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	dxxpdo_13;
input 	phi_mod_int_reg_8_3;
input 	dxxpdo_14;
input 	phi_mod_int_reg_9_3;
input 	dxxpdo_15;
input 	phi_mod_int_reg_10_3;
input 	dxxpdo_16;
input 	phi_mod_int_reg_11_3;
input 	dxxpdo_17;
input 	phi_mod_int_reg_12_3;
input 	dxxpdo_18;
input 	phi_mod_int_reg_13_3;
input 	dxxpdo_19;
input 	phi_mod_int_reg_14_3;
input 	dxxpdo_20;
input 	phi_mod_int_reg_15_3;
input 	dxxpdo_5;
input 	phi_mod_int_reg_0_3;
input 	dxxpdo_6;
input 	phi_mod_int_reg_1_3;
input 	dxxpdo_7;
input 	phi_mod_int_reg_2_3;
input 	dxxpdo_8;
input 	phi_mod_int_reg_3_3;
input 	dxxpdo_9;
input 	phi_mod_int_reg_4_3;
input 	dxxpdo_10;
input 	phi_mod_int_reg_5_3;
input 	dxxpdo_11;
input 	phi_mod_int_reg_6_3;
input 	dxxpdo_12;
input 	phi_mod_int_reg_7_3;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
input 	clock;
input 	clken;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~50 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~6 ;
wire \op_1~9_sumout ;
wire \op_1~10 ;
wire \op_1~13_sumout ;
wire \op_1~14 ;
wire \op_1~17_sumout ;
wire \op_1~18 ;
wire \op_1~21_sumout ;
wire \op_1~22 ;
wire \op_1~25_sumout ;
wire \op_1~26 ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;


dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_5),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_0_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_6),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_1_3),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_7),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_2_3),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_8),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_3_3),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_9),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_4_3),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

cyclonev_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_10),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_5_3),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

cyclonev_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_11),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_6_3),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

cyclonev_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_12),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_7_3),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_13),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_8_3),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_14),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_9_3),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_15),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_10_3),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_16),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_11_3),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_17),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_12_3),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_18),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_13_3),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_19),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_14_3),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_20),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_15_3),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

endmodule

module sine_mac_i_lpmd (
	q_a_0,
	q_b_0,
	q_a_1,
	q_b_1,
	q_a_2,
	q_b_2,
	q_a_3,
	q_b_3,
	q_a_4,
	q_b_4,
	q_a_5,
	q_b_5,
	q_a_6,
	q_b_6,
	q_a_7,
	q_b_7,
	q_a_8,
	q_b_8,
	q_a_9,
	q_b_9,
	q_a_10,
	q_b_10,
	q_a_11,
	q_b_11,
	q_a_12,
	q_b_12,
	q_a_13,
	q_b_13,
	q_a_14,
	q_b_14,
	q_a_15,
	q_b_15,
	q_a_16,
	q_b_16,
	q_a_17,
	q_b_17,
	q_a_18,
	q_b_18,
	q_a_19,
	q_b_19,
	q_a_20,
	q_b_20,
	q_a_21,
	q_b_21,
	q_a_22,
	q_b_22,
	q_a_23,
	q_b_23,
	q_a_01,
	q_a_110,
	q_a_24,
	q_a_31,
	q_a_41,
	q_a_51,
	q_a_61,
	q_a_71,
	q_a_81,
	q_a_91,
	q_a_101,
	q_a_111,
	q_a_121,
	q_a_131,
	q_a_141,
	q_a_151,
	q_a_161,
	q_a_171,
	q_a_181,
	q_a_191,
	q_a_201,
	q_a_211,
	q_a_221,
	q_a_231,
	q_a_02,
	q_a_112,
	q_a_25,
	q_a_32,
	q_a_42,
	q_a_52,
	q_a_62,
	q_a_72,
	q_a_82,
	q_a_92,
	q_a_102,
	q_a_113,
	q_a_122,
	q_a_132,
	q_a_142,
	q_a_152,
	q_a_162,
	q_a_172,
	q_a_182,
	q_a_192,
	q_a_202,
	q_a_212,
	q_a_222,
	q_a_232,
	dffe47,
	result_a_28,
	dffe24,
	dffe35,
	dffe48,
	dffe25,
	dffe26,
	dffe27,
	dffe28,
	dffe29,
	dffe30,
	dffe31,
	dffe32,
	dffe33,
	dffe34,
	dffe36,
	dffe37,
	dffe38,
	dffe39,
	dffe40,
	dffe41,
	dffe42,
	dffe43,
	dffe44,
	dffe45,
	dffe46,
	clk,
	clken,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	q_a_0;
input 	q_b_0;
input 	q_a_1;
input 	q_b_1;
input 	q_a_2;
input 	q_b_2;
input 	q_a_3;
input 	q_b_3;
input 	q_a_4;
input 	q_b_4;
input 	q_a_5;
input 	q_b_5;
input 	q_a_6;
input 	q_b_6;
input 	q_a_7;
input 	q_b_7;
input 	q_a_8;
input 	q_b_8;
input 	q_a_9;
input 	q_b_9;
input 	q_a_10;
input 	q_b_10;
input 	q_a_11;
input 	q_b_11;
input 	q_a_12;
input 	q_b_12;
input 	q_a_13;
input 	q_b_13;
input 	q_a_14;
input 	q_b_14;
input 	q_a_15;
input 	q_b_15;
input 	q_a_16;
input 	q_b_16;
input 	q_a_17;
input 	q_b_17;
input 	q_a_18;
input 	q_b_18;
input 	q_a_19;
input 	q_b_19;
input 	q_a_20;
input 	q_b_20;
input 	q_a_21;
input 	q_b_21;
input 	q_a_22;
input 	q_b_22;
input 	q_a_23;
input 	q_b_23;
input 	q_a_01;
input 	q_a_110;
input 	q_a_24;
input 	q_a_31;
input 	q_a_41;
input 	q_a_51;
input 	q_a_61;
input 	q_a_71;
input 	q_a_81;
input 	q_a_91;
input 	q_a_101;
input 	q_a_111;
input 	q_a_121;
input 	q_a_131;
input 	q_a_141;
input 	q_a_151;
input 	q_a_161;
input 	q_a_171;
input 	q_a_181;
input 	q_a_191;
input 	q_a_201;
input 	q_a_211;
input 	q_a_221;
input 	q_a_231;
input 	q_a_02;
input 	q_a_112;
input 	q_a_25;
input 	q_a_32;
input 	q_a_42;
input 	q_a_52;
input 	q_a_62;
input 	q_a_72;
input 	q_a_82;
input 	q_a_92;
input 	q_a_102;
input 	q_a_113;
input 	q_a_122;
input 	q_a_132;
input 	q_a_142;
input 	q_a_152;
input 	q_a_162;
input 	q_a_172;
input 	q_a_182;
input 	q_a_192;
input 	q_a_202;
input 	q_a_212;
input 	q_a_222;
input 	q_a_232;
output 	dffe47;
output 	result_a_28;
output 	dffe24;
output 	dffe35;
output 	dffe48;
output 	dffe25;
output 	dffe26;
output 	dffe27;
output 	dffe28;
output 	dffe29;
output 	dffe30;
output 	dffe31;
output 	dffe32;
output 	dffe33;
output 	dffe34;
output 	dffe36;
output 	dffe37;
output 	dffe38;
output 	dffe39;
output 	dffe40;
output 	dffe41;
output 	dffe42;
output 	dffe43;
output 	dffe44;
output 	dffe45;
output 	dffe46;
input 	clk;
input 	clken;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \result_a[46]~q ;
wire \result_b[46]~q ;
wire \result_a[23]~q ;
wire \result_b[23]~q ;
wire \result_a[34]~q ;
wire \result_b[34]~q ;
wire \result_a[47]~q ;
wire \result_b[47]~q ;
wire \result_a[24]~q ;
wire \result_b[24]~q ;
wire \result_a[25]~q ;
wire \result_b[25]~q ;
wire \result_a[26]~q ;
wire \result_b[26]~q ;
wire \result_a[27]~q ;
wire \result_b[27]~q ;
wire \result_a[28]~q ;
wire \result_b[28]~q ;
wire \result_a[29]~q ;
wire \result_b[29]~q ;
wire \result_a[30]~q ;
wire \result_b[30]~q ;
wire \result_a[31]~q ;
wire \result_b[31]~q ;
wire \result_a[32]~q ;
wire \result_b[32]~q ;
wire \result_a[33]~q ;
wire \result_b[33]~q ;
wire \result_a[35]~q ;
wire \result_b[35]~q ;
wire \result_a[36]~q ;
wire \result_b[36]~q ;
wire \result_a[37]~q ;
wire \result_b[37]~q ;
wire \result_a[38]~q ;
wire \result_b[38]~q ;
wire \result_a[39]~q ;
wire \result_b[39]~q ;
wire \result_a[40]~q ;
wire \result_b[40]~q ;
wire \result_a[41]~q ;
wire \result_b[41]~q ;
wire \result_a[42]~q ;
wire \result_b[42]~q ;
wire \result_a[43]~q ;
wire \result_b[43]~q ;
wire \result_a[44]~q ;
wire \result_b[44]~q ;
wire \result_a[45]~q ;
wire \result_b[45]~q ;
wire \result_a[22]~q ;
wire \result_b[22]~q ;
wire \result_a[21]~q ;
wire \result_b[21]~q ;
wire \result_a[20]~q ;
wire \result_b[20]~q ;
wire \result_a[19]~q ;
wire \result_b[19]~q ;
wire \result_a[18]~q ;
wire \result_b[18]~q ;
wire \result_a[17]~q ;
wire \result_b[17]~q ;
wire \result_a[16]~q ;
wire \result_b[16]~q ;
wire \result_a[15]~q ;
wire \result_b[15]~q ;
wire \result_a[14]~q ;
wire \result_b[14]~q ;
wire \result_a[13]~q ;
wire \result_b[13]~q ;
wire \result_a[12]~q ;
wire \result_b[12]~q ;
wire \result_a[11]~q ;
wire \result_b[11]~q ;
wire \result_a[10]~q ;
wire \result_b[10]~q ;
wire \result_a[9]~q ;
wire \result_b[9]~q ;
wire \result_a[8]~q ;
wire \result_b[8]~q ;
wire \result_a[7]~q ;
wire \result_b[7]~q ;
wire \result_a[6]~q ;
wire \result_b[6]~q ;
wire \result_a[5]~q ;
wire \result_b[5]~q ;
wire \result_a[4]~q ;
wire \result_b[4]~q ;
wire \result_a[3]~q ;
wire \result_b[3]~q ;
wire \result_a[2]~q ;
wire \result_b[2]~q ;
wire \result_a[1]~q ;
wire \result_b[1]~q ;
wire \result_a[0]~q ;
wire \result_b[0]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[46]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[46]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[23]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[23]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[34]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[34]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[47]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[47]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[24]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[24]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[25]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[25]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[26]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[26]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[27]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[27]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[28]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[28]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[29]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[29]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[30]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[30]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[31]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[31]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[32]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[32]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[33]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[33]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[35]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[35]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[36]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[36]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[37]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[37]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[38]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[38]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[39]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[39]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[40]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[40]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[41]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[41]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[42]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[42]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[43]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[43]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[44]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[44]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[45]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[45]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[22]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[22]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[21]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[21]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[20]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[20]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[19]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[19]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[18]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[18]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[17]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[17]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[16]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[16]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[15]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[15]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[14]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[14]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[13]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[13]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[12]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[12]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[11]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[11]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[10]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[10]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[9]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[9]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[8]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[8]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[7]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[7]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[6]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[6]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[5]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[5]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[4]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[4]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[3]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[3]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[2]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[2]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[1]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[1]~q ;
wire \m_0|lpm_mult_component|auto_generated|result_output_reg[0]~q ;
wire \m_1|lpm_mult_component|auto_generated|result_output_reg[0]~q ;


sine_las a_0(
	.result_a_46(\result_a[46]~q ),
	.result_b_46(\result_b[46]~q ),
	.result_a_23(\result_a[23]~q ),
	.result_b_23(\result_b[23]~q ),
	.result_a_34(\result_a[34]~q ),
	.result_b_34(\result_b[34]~q ),
	.result_a_47(\result_a[47]~q ),
	.result_b_47(\result_b[47]~q ),
	.result_a_24(\result_a[24]~q ),
	.result_b_24(\result_b[24]~q ),
	.result_a_25(\result_a[25]~q ),
	.result_b_25(\result_b[25]~q ),
	.result_a_26(\result_a[26]~q ),
	.result_b_26(\result_b[26]~q ),
	.result_a_27(\result_a[27]~q ),
	.result_b_27(\result_b[27]~q ),
	.result_a_28(\result_a[28]~q ),
	.result_b_28(\result_b[28]~q ),
	.result_a_29(\result_a[29]~q ),
	.result_b_29(\result_b[29]~q ),
	.result_a_30(\result_a[30]~q ),
	.result_b_30(\result_b[30]~q ),
	.result_a_31(\result_a[31]~q ),
	.result_b_31(\result_b[31]~q ),
	.result_a_32(\result_a[32]~q ),
	.result_b_32(\result_b[32]~q ),
	.result_a_33(\result_a[33]~q ),
	.result_b_33(\result_b[33]~q ),
	.result_a_35(\result_a[35]~q ),
	.result_b_35(\result_b[35]~q ),
	.result_a_36(\result_a[36]~q ),
	.result_b_36(\result_b[36]~q ),
	.result_a_37(\result_a[37]~q ),
	.result_b_37(\result_b[37]~q ),
	.result_a_38(\result_a[38]~q ),
	.result_b_38(\result_b[38]~q ),
	.result_a_39(\result_a[39]~q ),
	.result_b_39(\result_b[39]~q ),
	.result_a_40(\result_a[40]~q ),
	.result_b_40(\result_b[40]~q ),
	.result_a_41(\result_a[41]~q ),
	.result_b_41(\result_b[41]~q ),
	.result_a_42(\result_a[42]~q ),
	.result_b_42(\result_b[42]~q ),
	.result_a_43(\result_a[43]~q ),
	.result_b_43(\result_b[43]~q ),
	.result_a_44(\result_a[44]~q ),
	.result_b_44(\result_b[44]~q ),
	.result_a_45(\result_a[45]~q ),
	.result_b_45(\result_b[45]~q ),
	.result_a_22(\result_a[22]~q ),
	.result_b_22(\result_b[22]~q ),
	.result_a_21(\result_a[21]~q ),
	.result_b_21(\result_b[21]~q ),
	.result_a_20(\result_a[20]~q ),
	.result_b_20(\result_b[20]~q ),
	.result_a_19(\result_a[19]~q ),
	.result_b_19(\result_b[19]~q ),
	.result_a_18(\result_a[18]~q ),
	.result_b_18(\result_b[18]~q ),
	.result_a_17(\result_a[17]~q ),
	.result_b_17(\result_b[17]~q ),
	.result_a_16(\result_a[16]~q ),
	.result_b_16(\result_b[16]~q ),
	.result_a_15(\result_a[15]~q ),
	.result_b_15(\result_b[15]~q ),
	.result_a_14(\result_a[14]~q ),
	.result_b_14(\result_b[14]~q ),
	.result_a_13(\result_a[13]~q ),
	.result_b_13(\result_b[13]~q ),
	.result_a_12(\result_a[12]~q ),
	.result_b_12(\result_b[12]~q ),
	.result_a_11(\result_a[11]~q ),
	.result_b_11(\result_b[11]~q ),
	.result_a_10(\result_a[10]~q ),
	.result_b_10(\result_b[10]~q ),
	.result_a_9(\result_a[9]~q ),
	.result_b_9(\result_b[9]~q ),
	.result_a_8(\result_a[8]~q ),
	.result_b_8(\result_b[8]~q ),
	.result_a_7(\result_a[7]~q ),
	.result_b_7(\result_b[7]~q ),
	.result_a_6(\result_a[6]~q ),
	.result_b_6(\result_b[6]~q ),
	.result_a_5(\result_a[5]~q ),
	.result_b_5(\result_b[5]~q ),
	.result_a_4(\result_a[4]~q ),
	.result_b_4(\result_b[4]~q ),
	.result_a_3(\result_a[3]~q ),
	.result_b_3(\result_b[3]~q ),
	.result_a_2(\result_a[2]~q ),
	.result_b_2(\result_b[2]~q ),
	.result_a_1(\result_a[1]~q ),
	.result_b_1(\result_b[1]~q ),
	.result_a_0(\result_a[0]~q ),
	.result_b_0(\result_b[0]~q ),
	.dffe47(dffe47),
	.dffe24(dffe24),
	.dffe35(dffe35),
	.dffe48(dffe48),
	.dffe25(dffe25),
	.dffe26(dffe26),
	.dffe27(dffe27),
	.dffe28(dffe28),
	.dffe29(dffe29),
	.dffe30(dffe30),
	.dffe31(dffe31),
	.dffe32(dffe32),
	.dffe33(dffe33),
	.dffe34(dffe34),
	.dffe36(dffe36),
	.dffe37(dffe37),
	.dffe38(dffe38),
	.dffe39(dffe39),
	.dffe40(dffe40),
	.dffe41(dffe41),
	.dffe42(dffe42),
	.dffe43(dffe43),
	.dffe44(dffe44),
	.dffe45(dffe45),
	.dffe46(dffe46),
	.clk(clk),
	.clken(clken));

sine_lmsd_1 m_1(
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.q_b_22(q_b_22),
	.q_b_23(q_b_23),
	.q_a_0(q_a_02),
	.q_a_1(q_a_112),
	.q_a_2(q_a_25),
	.q_a_3(q_a_32),
	.q_a_4(q_a_42),
	.q_a_5(q_a_52),
	.q_a_6(q_a_62),
	.q_a_7(q_a_72),
	.q_a_8(q_a_82),
	.q_a_9(q_a_92),
	.q_a_10(q_a_102),
	.q_a_11(q_a_113),
	.q_a_12(q_a_122),
	.q_a_13(q_a_132),
	.q_a_14(q_a_142),
	.q_a_15(q_a_152),
	.q_a_16(q_a_162),
	.q_a_17(q_a_172),
	.q_a_18(q_a_182),
	.q_a_19(q_a_192),
	.q_a_20(q_a_202),
	.q_a_21(q_a_212),
	.q_a_22(q_a_222),
	.q_a_23(q_a_232),
	.result_output_reg_46(\m_1|lpm_mult_component|auto_generated|result_output_reg[46]~q ),
	.result_output_reg_23(\m_1|lpm_mult_component|auto_generated|result_output_reg[23]~q ),
	.result_output_reg_34(\m_1|lpm_mult_component|auto_generated|result_output_reg[34]~q ),
	.result_output_reg_47(\m_1|lpm_mult_component|auto_generated|result_output_reg[47]~q ),
	.result_output_reg_24(\m_1|lpm_mult_component|auto_generated|result_output_reg[24]~q ),
	.result_output_reg_25(\m_1|lpm_mult_component|auto_generated|result_output_reg[25]~q ),
	.result_output_reg_26(\m_1|lpm_mult_component|auto_generated|result_output_reg[26]~q ),
	.result_output_reg_27(\m_1|lpm_mult_component|auto_generated|result_output_reg[27]~q ),
	.result_output_reg_28(\m_1|lpm_mult_component|auto_generated|result_output_reg[28]~q ),
	.result_output_reg_29(\m_1|lpm_mult_component|auto_generated|result_output_reg[29]~q ),
	.result_output_reg_30(\m_1|lpm_mult_component|auto_generated|result_output_reg[30]~q ),
	.result_output_reg_31(\m_1|lpm_mult_component|auto_generated|result_output_reg[31]~q ),
	.result_output_reg_32(\m_1|lpm_mult_component|auto_generated|result_output_reg[32]~q ),
	.result_output_reg_33(\m_1|lpm_mult_component|auto_generated|result_output_reg[33]~q ),
	.result_output_reg_35(\m_1|lpm_mult_component|auto_generated|result_output_reg[35]~q ),
	.result_output_reg_36(\m_1|lpm_mult_component|auto_generated|result_output_reg[36]~q ),
	.result_output_reg_37(\m_1|lpm_mult_component|auto_generated|result_output_reg[37]~q ),
	.result_output_reg_38(\m_1|lpm_mult_component|auto_generated|result_output_reg[38]~q ),
	.result_output_reg_39(\m_1|lpm_mult_component|auto_generated|result_output_reg[39]~q ),
	.result_output_reg_40(\m_1|lpm_mult_component|auto_generated|result_output_reg[40]~q ),
	.result_output_reg_41(\m_1|lpm_mult_component|auto_generated|result_output_reg[41]~q ),
	.result_output_reg_42(\m_1|lpm_mult_component|auto_generated|result_output_reg[42]~q ),
	.result_output_reg_43(\m_1|lpm_mult_component|auto_generated|result_output_reg[43]~q ),
	.result_output_reg_44(\m_1|lpm_mult_component|auto_generated|result_output_reg[44]~q ),
	.result_output_reg_45(\m_1|lpm_mult_component|auto_generated|result_output_reg[45]~q ),
	.result_output_reg_22(\m_1|lpm_mult_component|auto_generated|result_output_reg[22]~q ),
	.result_output_reg_21(\m_1|lpm_mult_component|auto_generated|result_output_reg[21]~q ),
	.result_output_reg_20(\m_1|lpm_mult_component|auto_generated|result_output_reg[20]~q ),
	.result_output_reg_19(\m_1|lpm_mult_component|auto_generated|result_output_reg[19]~q ),
	.result_output_reg_18(\m_1|lpm_mult_component|auto_generated|result_output_reg[18]~q ),
	.result_output_reg_17(\m_1|lpm_mult_component|auto_generated|result_output_reg[17]~q ),
	.result_output_reg_16(\m_1|lpm_mult_component|auto_generated|result_output_reg[16]~q ),
	.result_output_reg_15(\m_1|lpm_mult_component|auto_generated|result_output_reg[15]~q ),
	.result_output_reg_14(\m_1|lpm_mult_component|auto_generated|result_output_reg[14]~q ),
	.result_output_reg_13(\m_1|lpm_mult_component|auto_generated|result_output_reg[13]~q ),
	.result_output_reg_12(\m_1|lpm_mult_component|auto_generated|result_output_reg[12]~q ),
	.result_output_reg_11(\m_1|lpm_mult_component|auto_generated|result_output_reg[11]~q ),
	.result_output_reg_10(\m_1|lpm_mult_component|auto_generated|result_output_reg[10]~q ),
	.result_output_reg_9(\m_1|lpm_mult_component|auto_generated|result_output_reg[9]~q ),
	.result_output_reg_8(\m_1|lpm_mult_component|auto_generated|result_output_reg[8]~q ),
	.result_output_reg_7(\m_1|lpm_mult_component|auto_generated|result_output_reg[7]~q ),
	.result_output_reg_6(\m_1|lpm_mult_component|auto_generated|result_output_reg[6]~q ),
	.result_output_reg_5(\m_1|lpm_mult_component|auto_generated|result_output_reg[5]~q ),
	.result_output_reg_4(\m_1|lpm_mult_component|auto_generated|result_output_reg[4]~q ),
	.result_output_reg_3(\m_1|lpm_mult_component|auto_generated|result_output_reg[3]~q ),
	.result_output_reg_2(\m_1|lpm_mult_component|auto_generated|result_output_reg[2]~q ),
	.result_output_reg_1(\m_1|lpm_mult_component|auto_generated|result_output_reg[1]~q ),
	.result_output_reg_0(\m_1|lpm_mult_component|auto_generated|result_output_reg[0]~q ),
	.clk(clk),
	.clken(clken));

sine_lmsd m_0(
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.q_a_8(q_a_8),
	.q_a_9(q_a_9),
	.q_a_10(q_a_10),
	.q_a_11(q_a_11),
	.q_a_12(q_a_12),
	.q_a_13(q_a_13),
	.q_a_14(q_a_14),
	.q_a_15(q_a_15),
	.q_a_16(q_a_16),
	.q_a_17(q_a_17),
	.q_a_18(q_a_18),
	.q_a_19(q_a_19),
	.q_a_20(q_a_20),
	.q_a_21(q_a_21),
	.q_a_22(q_a_22),
	.q_a_23(q_a_23),
	.q_a_01(q_a_01),
	.q_a_110(q_a_110),
	.q_a_24(q_a_24),
	.q_a_31(q_a_31),
	.q_a_41(q_a_41),
	.q_a_51(q_a_51),
	.q_a_61(q_a_61),
	.q_a_71(q_a_71),
	.q_a_81(q_a_81),
	.q_a_91(q_a_91),
	.q_a_101(q_a_101),
	.q_a_111(q_a_111),
	.q_a_121(q_a_121),
	.q_a_131(q_a_131),
	.q_a_141(q_a_141),
	.q_a_151(q_a_151),
	.q_a_161(q_a_161),
	.q_a_171(q_a_171),
	.q_a_181(q_a_181),
	.q_a_191(q_a_191),
	.q_a_201(q_a_201),
	.q_a_211(q_a_211),
	.q_a_221(q_a_221),
	.q_a_231(q_a_231),
	.result_output_reg_46(\m_0|lpm_mult_component|auto_generated|result_output_reg[46]~q ),
	.result_output_reg_23(\m_0|lpm_mult_component|auto_generated|result_output_reg[23]~q ),
	.result_output_reg_34(\m_0|lpm_mult_component|auto_generated|result_output_reg[34]~q ),
	.result_output_reg_47(\m_0|lpm_mult_component|auto_generated|result_output_reg[47]~q ),
	.result_output_reg_24(\m_0|lpm_mult_component|auto_generated|result_output_reg[24]~q ),
	.result_output_reg_25(\m_0|lpm_mult_component|auto_generated|result_output_reg[25]~q ),
	.result_output_reg_26(\m_0|lpm_mult_component|auto_generated|result_output_reg[26]~q ),
	.result_output_reg_27(\m_0|lpm_mult_component|auto_generated|result_output_reg[27]~q ),
	.result_output_reg_28(\m_0|lpm_mult_component|auto_generated|result_output_reg[28]~q ),
	.result_output_reg_29(\m_0|lpm_mult_component|auto_generated|result_output_reg[29]~q ),
	.result_output_reg_30(\m_0|lpm_mult_component|auto_generated|result_output_reg[30]~q ),
	.result_output_reg_31(\m_0|lpm_mult_component|auto_generated|result_output_reg[31]~q ),
	.result_output_reg_32(\m_0|lpm_mult_component|auto_generated|result_output_reg[32]~q ),
	.result_output_reg_33(\m_0|lpm_mult_component|auto_generated|result_output_reg[33]~q ),
	.result_output_reg_35(\m_0|lpm_mult_component|auto_generated|result_output_reg[35]~q ),
	.result_output_reg_36(\m_0|lpm_mult_component|auto_generated|result_output_reg[36]~q ),
	.result_output_reg_37(\m_0|lpm_mult_component|auto_generated|result_output_reg[37]~q ),
	.result_output_reg_38(\m_0|lpm_mult_component|auto_generated|result_output_reg[38]~q ),
	.result_output_reg_39(\m_0|lpm_mult_component|auto_generated|result_output_reg[39]~q ),
	.result_output_reg_40(\m_0|lpm_mult_component|auto_generated|result_output_reg[40]~q ),
	.result_output_reg_41(\m_0|lpm_mult_component|auto_generated|result_output_reg[41]~q ),
	.result_output_reg_42(\m_0|lpm_mult_component|auto_generated|result_output_reg[42]~q ),
	.result_output_reg_43(\m_0|lpm_mult_component|auto_generated|result_output_reg[43]~q ),
	.result_output_reg_44(\m_0|lpm_mult_component|auto_generated|result_output_reg[44]~q ),
	.result_output_reg_45(\m_0|lpm_mult_component|auto_generated|result_output_reg[45]~q ),
	.result_output_reg_22(\m_0|lpm_mult_component|auto_generated|result_output_reg[22]~q ),
	.result_output_reg_21(\m_0|lpm_mult_component|auto_generated|result_output_reg[21]~q ),
	.result_output_reg_20(\m_0|lpm_mult_component|auto_generated|result_output_reg[20]~q ),
	.result_output_reg_19(\m_0|lpm_mult_component|auto_generated|result_output_reg[19]~q ),
	.result_output_reg_18(\m_0|lpm_mult_component|auto_generated|result_output_reg[18]~q ),
	.result_output_reg_17(\m_0|lpm_mult_component|auto_generated|result_output_reg[17]~q ),
	.result_output_reg_16(\m_0|lpm_mult_component|auto_generated|result_output_reg[16]~q ),
	.result_output_reg_15(\m_0|lpm_mult_component|auto_generated|result_output_reg[15]~q ),
	.result_output_reg_14(\m_0|lpm_mult_component|auto_generated|result_output_reg[14]~q ),
	.result_output_reg_13(\m_0|lpm_mult_component|auto_generated|result_output_reg[13]~q ),
	.result_output_reg_12(\m_0|lpm_mult_component|auto_generated|result_output_reg[12]~q ),
	.result_output_reg_11(\m_0|lpm_mult_component|auto_generated|result_output_reg[11]~q ),
	.result_output_reg_10(\m_0|lpm_mult_component|auto_generated|result_output_reg[10]~q ),
	.result_output_reg_9(\m_0|lpm_mult_component|auto_generated|result_output_reg[9]~q ),
	.result_output_reg_8(\m_0|lpm_mult_component|auto_generated|result_output_reg[8]~q ),
	.result_output_reg_7(\m_0|lpm_mult_component|auto_generated|result_output_reg[7]~q ),
	.result_output_reg_6(\m_0|lpm_mult_component|auto_generated|result_output_reg[6]~q ),
	.result_output_reg_5(\m_0|lpm_mult_component|auto_generated|result_output_reg[5]~q ),
	.result_output_reg_4(\m_0|lpm_mult_component|auto_generated|result_output_reg[4]~q ),
	.result_output_reg_3(\m_0|lpm_mult_component|auto_generated|result_output_reg[3]~q ),
	.result_output_reg_2(\m_0|lpm_mult_component|auto_generated|result_output_reg[2]~q ),
	.result_output_reg_1(\m_0|lpm_mult_component|auto_generated|result_output_reg[1]~q ),
	.result_output_reg_0(\m_0|lpm_mult_component|auto_generated|result_output_reg[0]~q ),
	.clk(clk),
	.clken(clken));

dffeas \result_a[46] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[46]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[46]~q ),
	.prn(vcc));
defparam \result_a[46] .is_wysiwyg = "true";
defparam \result_a[46] .power_up = "low";

dffeas \result_b[46] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[46]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[46]~q ),
	.prn(vcc));
defparam \result_b[46] .is_wysiwyg = "true";
defparam \result_b[46] .power_up = "low";

dffeas \result_a[23] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[23]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[23]~q ),
	.prn(vcc));
defparam \result_a[23] .is_wysiwyg = "true";
defparam \result_a[23] .power_up = "low";

dffeas \result_b[23] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[23]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[23]~q ),
	.prn(vcc));
defparam \result_b[23] .is_wysiwyg = "true";
defparam \result_b[23] .power_up = "low";

dffeas \result_a[34] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[34]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[34]~q ),
	.prn(vcc));
defparam \result_a[34] .is_wysiwyg = "true";
defparam \result_a[34] .power_up = "low";

dffeas \result_b[34] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[34]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[34]~q ),
	.prn(vcc));
defparam \result_b[34] .is_wysiwyg = "true";
defparam \result_b[34] .power_up = "low";

dffeas \result_a[47] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[47]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[47]~q ),
	.prn(vcc));
defparam \result_a[47] .is_wysiwyg = "true";
defparam \result_a[47] .power_up = "low";

dffeas \result_b[47] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[47]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[47]~q ),
	.prn(vcc));
defparam \result_b[47] .is_wysiwyg = "true";
defparam \result_b[47] .power_up = "low";

dffeas \result_a[24] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[24]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[24]~q ),
	.prn(vcc));
defparam \result_a[24] .is_wysiwyg = "true";
defparam \result_a[24] .power_up = "low";

dffeas \result_b[24] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[24]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[24]~q ),
	.prn(vcc));
defparam \result_b[24] .is_wysiwyg = "true";
defparam \result_b[24] .power_up = "low";

dffeas \result_a[25] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[25]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[25]~q ),
	.prn(vcc));
defparam \result_a[25] .is_wysiwyg = "true";
defparam \result_a[25] .power_up = "low";

dffeas \result_b[25] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[25]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[25]~q ),
	.prn(vcc));
defparam \result_b[25] .is_wysiwyg = "true";
defparam \result_b[25] .power_up = "low";

dffeas \result_a[26] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[26]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[26]~q ),
	.prn(vcc));
defparam \result_a[26] .is_wysiwyg = "true";
defparam \result_a[26] .power_up = "low";

dffeas \result_b[26] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[26]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[26]~q ),
	.prn(vcc));
defparam \result_b[26] .is_wysiwyg = "true";
defparam \result_b[26] .power_up = "low";

dffeas \result_a[27] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[27]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[27]~q ),
	.prn(vcc));
defparam \result_a[27] .is_wysiwyg = "true";
defparam \result_a[27] .power_up = "low";

dffeas \result_b[27] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[27]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[27]~q ),
	.prn(vcc));
defparam \result_b[27] .is_wysiwyg = "true";
defparam \result_b[27] .power_up = "low";

dffeas \result_a[28] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[28]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[28]~q ),
	.prn(vcc));
defparam \result_a[28] .is_wysiwyg = "true";
defparam \result_a[28] .power_up = "low";

dffeas \result_b[28] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[28]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[28]~q ),
	.prn(vcc));
defparam \result_b[28] .is_wysiwyg = "true";
defparam \result_b[28] .power_up = "low";

dffeas \result_a[29] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[29]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[29]~q ),
	.prn(vcc));
defparam \result_a[29] .is_wysiwyg = "true";
defparam \result_a[29] .power_up = "low";

dffeas \result_b[29] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[29]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[29]~q ),
	.prn(vcc));
defparam \result_b[29] .is_wysiwyg = "true";
defparam \result_b[29] .power_up = "low";

dffeas \result_a[30] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[30]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[30]~q ),
	.prn(vcc));
defparam \result_a[30] .is_wysiwyg = "true";
defparam \result_a[30] .power_up = "low";

dffeas \result_b[30] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[30]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[30]~q ),
	.prn(vcc));
defparam \result_b[30] .is_wysiwyg = "true";
defparam \result_b[30] .power_up = "low";

dffeas \result_a[31] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[31]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[31]~q ),
	.prn(vcc));
defparam \result_a[31] .is_wysiwyg = "true";
defparam \result_a[31] .power_up = "low";

dffeas \result_b[31] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[31]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[31]~q ),
	.prn(vcc));
defparam \result_b[31] .is_wysiwyg = "true";
defparam \result_b[31] .power_up = "low";

dffeas \result_a[32] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[32]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[32]~q ),
	.prn(vcc));
defparam \result_a[32] .is_wysiwyg = "true";
defparam \result_a[32] .power_up = "low";

dffeas \result_b[32] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[32]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[32]~q ),
	.prn(vcc));
defparam \result_b[32] .is_wysiwyg = "true";
defparam \result_b[32] .power_up = "low";

dffeas \result_a[33] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[33]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[33]~q ),
	.prn(vcc));
defparam \result_a[33] .is_wysiwyg = "true";
defparam \result_a[33] .power_up = "low";

dffeas \result_b[33] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[33]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[33]~q ),
	.prn(vcc));
defparam \result_b[33] .is_wysiwyg = "true";
defparam \result_b[33] .power_up = "low";

dffeas \result_a[35] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[35]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[35]~q ),
	.prn(vcc));
defparam \result_a[35] .is_wysiwyg = "true";
defparam \result_a[35] .power_up = "low";

dffeas \result_b[35] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[35]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[35]~q ),
	.prn(vcc));
defparam \result_b[35] .is_wysiwyg = "true";
defparam \result_b[35] .power_up = "low";

dffeas \result_a[36] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[36]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[36]~q ),
	.prn(vcc));
defparam \result_a[36] .is_wysiwyg = "true";
defparam \result_a[36] .power_up = "low";

dffeas \result_b[36] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[36]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[36]~q ),
	.prn(vcc));
defparam \result_b[36] .is_wysiwyg = "true";
defparam \result_b[36] .power_up = "low";

dffeas \result_a[37] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[37]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[37]~q ),
	.prn(vcc));
defparam \result_a[37] .is_wysiwyg = "true";
defparam \result_a[37] .power_up = "low";

dffeas \result_b[37] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[37]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[37]~q ),
	.prn(vcc));
defparam \result_b[37] .is_wysiwyg = "true";
defparam \result_b[37] .power_up = "low";

dffeas \result_a[38] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[38]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[38]~q ),
	.prn(vcc));
defparam \result_a[38] .is_wysiwyg = "true";
defparam \result_a[38] .power_up = "low";

dffeas \result_b[38] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[38]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[38]~q ),
	.prn(vcc));
defparam \result_b[38] .is_wysiwyg = "true";
defparam \result_b[38] .power_up = "low";

dffeas \result_a[39] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[39]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[39]~q ),
	.prn(vcc));
defparam \result_a[39] .is_wysiwyg = "true";
defparam \result_a[39] .power_up = "low";

dffeas \result_b[39] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[39]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[39]~q ),
	.prn(vcc));
defparam \result_b[39] .is_wysiwyg = "true";
defparam \result_b[39] .power_up = "low";

dffeas \result_a[40] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[40]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[40]~q ),
	.prn(vcc));
defparam \result_a[40] .is_wysiwyg = "true";
defparam \result_a[40] .power_up = "low";

dffeas \result_b[40] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[40]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[40]~q ),
	.prn(vcc));
defparam \result_b[40] .is_wysiwyg = "true";
defparam \result_b[40] .power_up = "low";

dffeas \result_a[41] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[41]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[41]~q ),
	.prn(vcc));
defparam \result_a[41] .is_wysiwyg = "true";
defparam \result_a[41] .power_up = "low";

dffeas \result_b[41] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[41]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[41]~q ),
	.prn(vcc));
defparam \result_b[41] .is_wysiwyg = "true";
defparam \result_b[41] .power_up = "low";

dffeas \result_a[42] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[42]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[42]~q ),
	.prn(vcc));
defparam \result_a[42] .is_wysiwyg = "true";
defparam \result_a[42] .power_up = "low";

dffeas \result_b[42] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[42]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[42]~q ),
	.prn(vcc));
defparam \result_b[42] .is_wysiwyg = "true";
defparam \result_b[42] .power_up = "low";

dffeas \result_a[43] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[43]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[43]~q ),
	.prn(vcc));
defparam \result_a[43] .is_wysiwyg = "true";
defparam \result_a[43] .power_up = "low";

dffeas \result_b[43] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[43]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[43]~q ),
	.prn(vcc));
defparam \result_b[43] .is_wysiwyg = "true";
defparam \result_b[43] .power_up = "low";

dffeas \result_a[44] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[44]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[44]~q ),
	.prn(vcc));
defparam \result_a[44] .is_wysiwyg = "true";
defparam \result_a[44] .power_up = "low";

dffeas \result_b[44] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[44]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[44]~q ),
	.prn(vcc));
defparam \result_b[44] .is_wysiwyg = "true";
defparam \result_b[44] .power_up = "low";

dffeas \result_a[45] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[45]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[45]~q ),
	.prn(vcc));
defparam \result_a[45] .is_wysiwyg = "true";
defparam \result_a[45] .power_up = "low";

dffeas \result_b[45] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[45]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[45]~q ),
	.prn(vcc));
defparam \result_b[45] .is_wysiwyg = "true";
defparam \result_b[45] .power_up = "low";

dffeas \result_a[22] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[22]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[22]~q ),
	.prn(vcc));
defparam \result_a[22] .is_wysiwyg = "true";
defparam \result_a[22] .power_up = "low";

dffeas \result_b[22] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[22]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[22]~q ),
	.prn(vcc));
defparam \result_b[22] .is_wysiwyg = "true";
defparam \result_b[22] .power_up = "low";

dffeas \result_a[21] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[21]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[21]~q ),
	.prn(vcc));
defparam \result_a[21] .is_wysiwyg = "true";
defparam \result_a[21] .power_up = "low";

dffeas \result_b[21] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[21]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[21]~q ),
	.prn(vcc));
defparam \result_b[21] .is_wysiwyg = "true";
defparam \result_b[21] .power_up = "low";

dffeas \result_a[20] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[20]~q ),
	.prn(vcc));
defparam \result_a[20] .is_wysiwyg = "true";
defparam \result_a[20] .power_up = "low";

dffeas \result_b[20] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[20]~q ),
	.prn(vcc));
defparam \result_b[20] .is_wysiwyg = "true";
defparam \result_b[20] .power_up = "low";

dffeas \result_a[19] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[19]~q ),
	.prn(vcc));
defparam \result_a[19] .is_wysiwyg = "true";
defparam \result_a[19] .power_up = "low";

dffeas \result_b[19] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[19]~q ),
	.prn(vcc));
defparam \result_b[19] .is_wysiwyg = "true";
defparam \result_b[19] .power_up = "low";

dffeas \result_a[18] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[18]~q ),
	.prn(vcc));
defparam \result_a[18] .is_wysiwyg = "true";
defparam \result_a[18] .power_up = "low";

dffeas \result_b[18] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[18]~q ),
	.prn(vcc));
defparam \result_b[18] .is_wysiwyg = "true";
defparam \result_b[18] .power_up = "low";

dffeas \result_a[17] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[17]~q ),
	.prn(vcc));
defparam \result_a[17] .is_wysiwyg = "true";
defparam \result_a[17] .power_up = "low";

dffeas \result_b[17] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[17]~q ),
	.prn(vcc));
defparam \result_b[17] .is_wysiwyg = "true";
defparam \result_b[17] .power_up = "low";

dffeas \result_a[16] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[16]~q ),
	.prn(vcc));
defparam \result_a[16] .is_wysiwyg = "true";
defparam \result_a[16] .power_up = "low";

dffeas \result_b[16] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[16]~q ),
	.prn(vcc));
defparam \result_b[16] .is_wysiwyg = "true";
defparam \result_b[16] .power_up = "low";

dffeas \result_a[15] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[15]~q ),
	.prn(vcc));
defparam \result_a[15] .is_wysiwyg = "true";
defparam \result_a[15] .power_up = "low";

dffeas \result_b[15] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[15]~q ),
	.prn(vcc));
defparam \result_b[15] .is_wysiwyg = "true";
defparam \result_b[15] .power_up = "low";

dffeas \result_a[14] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[14]~q ),
	.prn(vcc));
defparam \result_a[14] .is_wysiwyg = "true";
defparam \result_a[14] .power_up = "low";

dffeas \result_b[14] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[14]~q ),
	.prn(vcc));
defparam \result_b[14] .is_wysiwyg = "true";
defparam \result_b[14] .power_up = "low";

dffeas \result_a[13] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[13]~q ),
	.prn(vcc));
defparam \result_a[13] .is_wysiwyg = "true";
defparam \result_a[13] .power_up = "low";

dffeas \result_b[13] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[13]~q ),
	.prn(vcc));
defparam \result_b[13] .is_wysiwyg = "true";
defparam \result_b[13] .power_up = "low";

dffeas \result_a[12] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[12]~q ),
	.prn(vcc));
defparam \result_a[12] .is_wysiwyg = "true";
defparam \result_a[12] .power_up = "low";

dffeas \result_b[12] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[12]~q ),
	.prn(vcc));
defparam \result_b[12] .is_wysiwyg = "true";
defparam \result_b[12] .power_up = "low";

dffeas \result_a[11] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[11]~q ),
	.prn(vcc));
defparam \result_a[11] .is_wysiwyg = "true";
defparam \result_a[11] .power_up = "low";

dffeas \result_b[11] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[11]~q ),
	.prn(vcc));
defparam \result_b[11] .is_wysiwyg = "true";
defparam \result_b[11] .power_up = "low";

dffeas \result_a[10] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[10]~q ),
	.prn(vcc));
defparam \result_a[10] .is_wysiwyg = "true";
defparam \result_a[10] .power_up = "low";

dffeas \result_b[10] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[10]~q ),
	.prn(vcc));
defparam \result_b[10] .is_wysiwyg = "true";
defparam \result_b[10] .power_up = "low";

dffeas \result_a[9] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[9]~q ),
	.prn(vcc));
defparam \result_a[9] .is_wysiwyg = "true";
defparam \result_a[9] .power_up = "low";

dffeas \result_b[9] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[9]~q ),
	.prn(vcc));
defparam \result_b[9] .is_wysiwyg = "true";
defparam \result_b[9] .power_up = "low";

dffeas \result_a[8] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[8]~q ),
	.prn(vcc));
defparam \result_a[8] .is_wysiwyg = "true";
defparam \result_a[8] .power_up = "low";

dffeas \result_b[8] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[8]~q ),
	.prn(vcc));
defparam \result_b[8] .is_wysiwyg = "true";
defparam \result_b[8] .power_up = "low";

dffeas \result_a[7] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[7]~q ),
	.prn(vcc));
defparam \result_a[7] .is_wysiwyg = "true";
defparam \result_a[7] .power_up = "low";

dffeas \result_b[7] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[7]~q ),
	.prn(vcc));
defparam \result_b[7] .is_wysiwyg = "true";
defparam \result_b[7] .power_up = "low";

dffeas \result_a[6] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[6]~q ),
	.prn(vcc));
defparam \result_a[6] .is_wysiwyg = "true";
defparam \result_a[6] .power_up = "low";

dffeas \result_b[6] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[6]~q ),
	.prn(vcc));
defparam \result_b[6] .is_wysiwyg = "true";
defparam \result_b[6] .power_up = "low";

dffeas \result_a[5] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[5]~q ),
	.prn(vcc));
defparam \result_a[5] .is_wysiwyg = "true";
defparam \result_a[5] .power_up = "low";

dffeas \result_b[5] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[5]~q ),
	.prn(vcc));
defparam \result_b[5] .is_wysiwyg = "true";
defparam \result_b[5] .power_up = "low";

dffeas \result_a[4] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[4]~q ),
	.prn(vcc));
defparam \result_a[4] .is_wysiwyg = "true";
defparam \result_a[4] .power_up = "low";

dffeas \result_b[4] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[4]~q ),
	.prn(vcc));
defparam \result_b[4] .is_wysiwyg = "true";
defparam \result_b[4] .power_up = "low";

dffeas \result_a[3] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[3]~q ),
	.prn(vcc));
defparam \result_a[3] .is_wysiwyg = "true";
defparam \result_a[3] .power_up = "low";

dffeas \result_b[3] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[3]~q ),
	.prn(vcc));
defparam \result_b[3] .is_wysiwyg = "true";
defparam \result_b[3] .power_up = "low";

dffeas \result_a[2] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[2]~q ),
	.prn(vcc));
defparam \result_a[2] .is_wysiwyg = "true";
defparam \result_a[2] .power_up = "low";

dffeas \result_b[2] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[2]~q ),
	.prn(vcc));
defparam \result_b[2] .is_wysiwyg = "true";
defparam \result_b[2] .power_up = "low";

dffeas \result_a[1] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[1]~q ),
	.prn(vcc));
defparam \result_a[1] .is_wysiwyg = "true";
defparam \result_a[1] .power_up = "low";

dffeas \result_b[1] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[1]~q ),
	.prn(vcc));
defparam \result_b[1] .is_wysiwyg = "true";
defparam \result_b[1] .power_up = "low";

dffeas \result_a[0] (
	.clk(clk),
	.d(\m_0|lpm_mult_component|auto_generated|result_output_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_a[0]~q ),
	.prn(vcc));
defparam \result_a[0] .is_wysiwyg = "true";
defparam \result_a[0] .power_up = "low";

dffeas \result_b[0] (
	.clk(clk),
	.d(\m_1|lpm_mult_component|auto_generated|result_output_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(result_a_28),
	.q(\result_b[0]~q ),
	.prn(vcc));
defparam \result_b[0] .is_wysiwyg = "true";
defparam \result_b[0] .power_up = "low";

cyclonev_lcell_comb \result_a[28]~0 (
	.dataa(!clken),
	.datab(!reset_n),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(result_a_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \result_a[28]~0 .extended_lut = "off";
defparam \result_a[28]~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \result_a[28]~0 .shared_arith = "off";

endmodule

module sine_las (
	result_a_46,
	result_b_46,
	result_a_23,
	result_b_23,
	result_a_34,
	result_b_34,
	result_a_47,
	result_b_47,
	result_a_24,
	result_b_24,
	result_a_25,
	result_b_25,
	result_a_26,
	result_b_26,
	result_a_27,
	result_b_27,
	result_a_28,
	result_b_28,
	result_a_29,
	result_b_29,
	result_a_30,
	result_b_30,
	result_a_31,
	result_b_31,
	result_a_32,
	result_b_32,
	result_a_33,
	result_b_33,
	result_a_35,
	result_b_35,
	result_a_36,
	result_b_36,
	result_a_37,
	result_b_37,
	result_a_38,
	result_b_38,
	result_a_39,
	result_b_39,
	result_a_40,
	result_b_40,
	result_a_41,
	result_b_41,
	result_a_42,
	result_b_42,
	result_a_43,
	result_b_43,
	result_a_44,
	result_b_44,
	result_a_45,
	result_b_45,
	result_a_22,
	result_b_22,
	result_a_21,
	result_b_21,
	result_a_20,
	result_b_20,
	result_a_19,
	result_b_19,
	result_a_18,
	result_b_18,
	result_a_17,
	result_b_17,
	result_a_16,
	result_b_16,
	result_a_15,
	result_b_15,
	result_a_14,
	result_b_14,
	result_a_13,
	result_b_13,
	result_a_12,
	result_b_12,
	result_a_11,
	result_b_11,
	result_a_10,
	result_b_10,
	result_a_9,
	result_b_9,
	result_a_8,
	result_b_8,
	result_a_7,
	result_b_7,
	result_a_6,
	result_b_6,
	result_a_5,
	result_b_5,
	result_a_4,
	result_b_4,
	result_a_3,
	result_b_3,
	result_a_2,
	result_b_2,
	result_a_1,
	result_b_1,
	result_a_0,
	result_b_0,
	dffe47,
	dffe24,
	dffe35,
	dffe48,
	dffe25,
	dffe26,
	dffe27,
	dffe28,
	dffe29,
	dffe30,
	dffe31,
	dffe32,
	dffe33,
	dffe34,
	dffe36,
	dffe37,
	dffe38,
	dffe39,
	dffe40,
	dffe41,
	dffe42,
	dffe43,
	dffe44,
	dffe45,
	dffe46,
	clk,
	clken)/* synthesis synthesis_greybox=1 */;
input 	result_a_46;
input 	result_b_46;
input 	result_a_23;
input 	result_b_23;
input 	result_a_34;
input 	result_b_34;
input 	result_a_47;
input 	result_b_47;
input 	result_a_24;
input 	result_b_24;
input 	result_a_25;
input 	result_b_25;
input 	result_a_26;
input 	result_b_26;
input 	result_a_27;
input 	result_b_27;
input 	result_a_28;
input 	result_b_28;
input 	result_a_29;
input 	result_b_29;
input 	result_a_30;
input 	result_b_30;
input 	result_a_31;
input 	result_b_31;
input 	result_a_32;
input 	result_b_32;
input 	result_a_33;
input 	result_b_33;
input 	result_a_35;
input 	result_b_35;
input 	result_a_36;
input 	result_b_36;
input 	result_a_37;
input 	result_b_37;
input 	result_a_38;
input 	result_b_38;
input 	result_a_39;
input 	result_b_39;
input 	result_a_40;
input 	result_b_40;
input 	result_a_41;
input 	result_b_41;
input 	result_a_42;
input 	result_b_42;
input 	result_a_43;
input 	result_b_43;
input 	result_a_44;
input 	result_b_44;
input 	result_a_45;
input 	result_b_45;
input 	result_a_22;
input 	result_b_22;
input 	result_a_21;
input 	result_b_21;
input 	result_a_20;
input 	result_b_20;
input 	result_a_19;
input 	result_b_19;
input 	result_a_18;
input 	result_b_18;
input 	result_a_17;
input 	result_b_17;
input 	result_a_16;
input 	result_b_16;
input 	result_a_15;
input 	result_b_15;
input 	result_a_14;
input 	result_b_14;
input 	result_a_13;
input 	result_b_13;
input 	result_a_12;
input 	result_b_12;
input 	result_a_11;
input 	result_b_11;
input 	result_a_10;
input 	result_b_10;
input 	result_a_9;
input 	result_b_9;
input 	result_a_8;
input 	result_b_8;
input 	result_a_7;
input 	result_b_7;
input 	result_a_6;
input 	result_b_6;
input 	result_a_5;
input 	result_b_5;
input 	result_a_4;
input 	result_b_4;
input 	result_a_3;
input 	result_b_3;
input 	result_a_2;
input 	result_b_2;
input 	result_a_1;
input 	result_b_1;
input 	result_a_0;
input 	result_b_0;
output 	dffe47;
output 	dffe24;
output 	dffe35;
output 	dffe48;
output 	dffe25;
output 	dffe26;
output 	dffe27;
output 	dffe28;
output 	dffe29;
output 	dffe30;
output 	dffe31;
output 	dffe32;
output 	dffe33;
output 	dffe34;
output 	dffe36;
output 	dffe37;
output 	dffe38;
output 	dffe39;
output 	dffe40;
output 	dffe41;
output 	dffe42;
output 	dffe43;
output 	dffe44;
output 	dffe45;
output 	dffe46;
input 	clk;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_lpm_add_sub_5 lpm_add_sub_component(
	.result_a_46(result_a_46),
	.result_b_46(result_b_46),
	.result_a_23(result_a_23),
	.result_b_23(result_b_23),
	.result_a_34(result_a_34),
	.result_b_34(result_b_34),
	.result_a_47(result_a_47),
	.result_b_47(result_b_47),
	.result_a_24(result_a_24),
	.result_b_24(result_b_24),
	.result_a_25(result_a_25),
	.result_b_25(result_b_25),
	.result_a_26(result_a_26),
	.result_b_26(result_b_26),
	.result_a_27(result_a_27),
	.result_b_27(result_b_27),
	.result_a_28(result_a_28),
	.result_b_28(result_b_28),
	.result_a_29(result_a_29),
	.result_b_29(result_b_29),
	.result_a_30(result_a_30),
	.result_b_30(result_b_30),
	.result_a_31(result_a_31),
	.result_b_31(result_b_31),
	.result_a_32(result_a_32),
	.result_b_32(result_b_32),
	.result_a_33(result_a_33),
	.result_b_33(result_b_33),
	.result_a_35(result_a_35),
	.result_b_35(result_b_35),
	.result_a_36(result_a_36),
	.result_b_36(result_b_36),
	.result_a_37(result_a_37),
	.result_b_37(result_b_37),
	.result_a_38(result_a_38),
	.result_b_38(result_b_38),
	.result_a_39(result_a_39),
	.result_b_39(result_b_39),
	.result_a_40(result_a_40),
	.result_b_40(result_b_40),
	.result_a_41(result_a_41),
	.result_b_41(result_b_41),
	.result_a_42(result_a_42),
	.result_b_42(result_b_42),
	.result_a_43(result_a_43),
	.result_b_43(result_b_43),
	.result_a_44(result_a_44),
	.result_b_44(result_b_44),
	.result_a_45(result_a_45),
	.result_b_45(result_b_45),
	.result_a_22(result_a_22),
	.result_b_22(result_b_22),
	.result_a_21(result_a_21),
	.result_b_21(result_b_21),
	.result_a_20(result_a_20),
	.result_b_20(result_b_20),
	.result_a_19(result_a_19),
	.result_b_19(result_b_19),
	.result_a_18(result_a_18),
	.result_b_18(result_b_18),
	.result_a_17(result_a_17),
	.result_b_17(result_b_17),
	.result_a_16(result_a_16),
	.result_b_16(result_b_16),
	.result_a_15(result_a_15),
	.result_b_15(result_b_15),
	.result_a_14(result_a_14),
	.result_b_14(result_b_14),
	.result_a_13(result_a_13),
	.result_b_13(result_b_13),
	.result_a_12(result_a_12),
	.result_b_12(result_b_12),
	.result_a_11(result_a_11),
	.result_b_11(result_b_11),
	.result_a_10(result_a_10),
	.result_b_10(result_b_10),
	.result_a_9(result_a_9),
	.result_b_9(result_b_9),
	.result_a_8(result_a_8),
	.result_b_8(result_b_8),
	.result_a_7(result_a_7),
	.result_b_7(result_b_7),
	.result_a_6(result_a_6),
	.result_b_6(result_b_6),
	.result_a_5(result_a_5),
	.result_b_5(result_b_5),
	.result_a_4(result_a_4),
	.result_b_4(result_b_4),
	.result_a_3(result_a_3),
	.result_b_3(result_b_3),
	.result_a_2(result_a_2),
	.result_b_2(result_b_2),
	.result_a_1(result_a_1),
	.result_b_1(result_b_1),
	.result_a_0(result_a_0),
	.result_b_0(result_b_0),
	.dffe47(dffe47),
	.dffe24(dffe24),
	.dffe35(dffe35),
	.dffe48(dffe48),
	.dffe25(dffe25),
	.dffe26(dffe26),
	.dffe27(dffe27),
	.dffe28(dffe28),
	.dffe29(dffe29),
	.dffe30(dffe30),
	.dffe31(dffe31),
	.dffe32(dffe32),
	.dffe33(dffe33),
	.dffe34(dffe34),
	.dffe36(dffe36),
	.dffe37(dffe37),
	.dffe38(dffe38),
	.dffe39(dffe39),
	.dffe40(dffe40),
	.dffe41(dffe41),
	.dffe42(dffe42),
	.dffe43(dffe43),
	.dffe44(dffe44),
	.dffe45(dffe45),
	.dffe46(dffe46),
	.clock(clk),
	.clken(clken));

endmodule

module sine_lpm_add_sub_5 (
	result_a_46,
	result_b_46,
	result_a_23,
	result_b_23,
	result_a_34,
	result_b_34,
	result_a_47,
	result_b_47,
	result_a_24,
	result_b_24,
	result_a_25,
	result_b_25,
	result_a_26,
	result_b_26,
	result_a_27,
	result_b_27,
	result_a_28,
	result_b_28,
	result_a_29,
	result_b_29,
	result_a_30,
	result_b_30,
	result_a_31,
	result_b_31,
	result_a_32,
	result_b_32,
	result_a_33,
	result_b_33,
	result_a_35,
	result_b_35,
	result_a_36,
	result_b_36,
	result_a_37,
	result_b_37,
	result_a_38,
	result_b_38,
	result_a_39,
	result_b_39,
	result_a_40,
	result_b_40,
	result_a_41,
	result_b_41,
	result_a_42,
	result_b_42,
	result_a_43,
	result_b_43,
	result_a_44,
	result_b_44,
	result_a_45,
	result_b_45,
	result_a_22,
	result_b_22,
	result_a_21,
	result_b_21,
	result_a_20,
	result_b_20,
	result_a_19,
	result_b_19,
	result_a_18,
	result_b_18,
	result_a_17,
	result_b_17,
	result_a_16,
	result_b_16,
	result_a_15,
	result_b_15,
	result_a_14,
	result_b_14,
	result_a_13,
	result_b_13,
	result_a_12,
	result_b_12,
	result_a_11,
	result_b_11,
	result_a_10,
	result_b_10,
	result_a_9,
	result_b_9,
	result_a_8,
	result_b_8,
	result_a_7,
	result_b_7,
	result_a_6,
	result_b_6,
	result_a_5,
	result_b_5,
	result_a_4,
	result_b_4,
	result_a_3,
	result_b_3,
	result_a_2,
	result_b_2,
	result_a_1,
	result_b_1,
	result_a_0,
	result_b_0,
	dffe47,
	dffe24,
	dffe35,
	dffe48,
	dffe25,
	dffe26,
	dffe27,
	dffe28,
	dffe29,
	dffe30,
	dffe31,
	dffe32,
	dffe33,
	dffe34,
	dffe36,
	dffe37,
	dffe38,
	dffe39,
	dffe40,
	dffe41,
	dffe42,
	dffe43,
	dffe44,
	dffe45,
	dffe46,
	clock,
	clken)/* synthesis synthesis_greybox=1 */;
input 	result_a_46;
input 	result_b_46;
input 	result_a_23;
input 	result_b_23;
input 	result_a_34;
input 	result_b_34;
input 	result_a_47;
input 	result_b_47;
input 	result_a_24;
input 	result_b_24;
input 	result_a_25;
input 	result_b_25;
input 	result_a_26;
input 	result_b_26;
input 	result_a_27;
input 	result_b_27;
input 	result_a_28;
input 	result_b_28;
input 	result_a_29;
input 	result_b_29;
input 	result_a_30;
input 	result_b_30;
input 	result_a_31;
input 	result_b_31;
input 	result_a_32;
input 	result_b_32;
input 	result_a_33;
input 	result_b_33;
input 	result_a_35;
input 	result_b_35;
input 	result_a_36;
input 	result_b_36;
input 	result_a_37;
input 	result_b_37;
input 	result_a_38;
input 	result_b_38;
input 	result_a_39;
input 	result_b_39;
input 	result_a_40;
input 	result_b_40;
input 	result_a_41;
input 	result_b_41;
input 	result_a_42;
input 	result_b_42;
input 	result_a_43;
input 	result_b_43;
input 	result_a_44;
input 	result_b_44;
input 	result_a_45;
input 	result_b_45;
input 	result_a_22;
input 	result_b_22;
input 	result_a_21;
input 	result_b_21;
input 	result_a_20;
input 	result_b_20;
input 	result_a_19;
input 	result_b_19;
input 	result_a_18;
input 	result_b_18;
input 	result_a_17;
input 	result_b_17;
input 	result_a_16;
input 	result_b_16;
input 	result_a_15;
input 	result_b_15;
input 	result_a_14;
input 	result_b_14;
input 	result_a_13;
input 	result_b_13;
input 	result_a_12;
input 	result_b_12;
input 	result_a_11;
input 	result_b_11;
input 	result_a_10;
input 	result_b_10;
input 	result_a_9;
input 	result_b_9;
input 	result_a_8;
input 	result_b_8;
input 	result_a_7;
input 	result_b_7;
input 	result_a_6;
input 	result_b_6;
input 	result_a_5;
input 	result_b_5;
input 	result_a_4;
input 	result_b_4;
input 	result_a_3;
input 	result_b_3;
input 	result_a_2;
input 	result_b_2;
input 	result_a_1;
input 	result_b_1;
input 	result_a_0;
input 	result_b_0;
output 	dffe47;
output 	dffe24;
output 	dffe35;
output 	dffe48;
output 	dffe25;
output 	dffe26;
output 	dffe27;
output 	dffe28;
output 	dffe29;
output 	dffe30;
output 	dffe31;
output 	dffe32;
output 	dffe33;
output 	dffe34;
output 	dffe36;
output 	dffe37;
output 	dffe38;
output 	dffe39;
output 	dffe40;
output 	dffe41;
output 	dffe42;
output 	dffe43;
output 	dffe44;
output 	dffe45;
output 	dffe46;
input 	clock;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_add_sub_5pi auto_generated(
	.result_a_46(result_a_46),
	.result_b_46(result_b_46),
	.result_a_23(result_a_23),
	.result_b_23(result_b_23),
	.result_a_34(result_a_34),
	.result_b_34(result_b_34),
	.result_a_47(result_a_47),
	.result_b_47(result_b_47),
	.result_a_24(result_a_24),
	.result_b_24(result_b_24),
	.result_a_25(result_a_25),
	.result_b_25(result_b_25),
	.result_a_26(result_a_26),
	.result_b_26(result_b_26),
	.result_a_27(result_a_27),
	.result_b_27(result_b_27),
	.result_a_28(result_a_28),
	.result_b_28(result_b_28),
	.result_a_29(result_a_29),
	.result_b_29(result_b_29),
	.result_a_30(result_a_30),
	.result_b_30(result_b_30),
	.result_a_31(result_a_31),
	.result_b_31(result_b_31),
	.result_a_32(result_a_32),
	.result_b_32(result_b_32),
	.result_a_33(result_a_33),
	.result_b_33(result_b_33),
	.result_a_35(result_a_35),
	.result_b_35(result_b_35),
	.result_a_36(result_a_36),
	.result_b_36(result_b_36),
	.result_a_37(result_a_37),
	.result_b_37(result_b_37),
	.result_a_38(result_a_38),
	.result_b_38(result_b_38),
	.result_a_39(result_a_39),
	.result_b_39(result_b_39),
	.result_a_40(result_a_40),
	.result_b_40(result_b_40),
	.result_a_41(result_a_41),
	.result_b_41(result_b_41),
	.result_a_42(result_a_42),
	.result_b_42(result_b_42),
	.result_a_43(result_a_43),
	.result_b_43(result_b_43),
	.result_a_44(result_a_44),
	.result_b_44(result_b_44),
	.result_a_45(result_a_45),
	.result_b_45(result_b_45),
	.result_a_22(result_a_22),
	.result_b_22(result_b_22),
	.result_a_21(result_a_21),
	.result_b_21(result_b_21),
	.result_a_20(result_a_20),
	.result_b_20(result_b_20),
	.result_a_19(result_a_19),
	.result_b_19(result_b_19),
	.result_a_18(result_a_18),
	.result_b_18(result_b_18),
	.result_a_17(result_a_17),
	.result_b_17(result_b_17),
	.result_a_16(result_a_16),
	.result_b_16(result_b_16),
	.result_a_15(result_a_15),
	.result_b_15(result_b_15),
	.result_a_14(result_a_14),
	.result_b_14(result_b_14),
	.result_a_13(result_a_13),
	.result_b_13(result_b_13),
	.result_a_12(result_a_12),
	.result_b_12(result_b_12),
	.result_a_11(result_a_11),
	.result_b_11(result_b_11),
	.result_a_10(result_a_10),
	.result_b_10(result_b_10),
	.result_a_9(result_a_9),
	.result_b_9(result_b_9),
	.result_a_8(result_a_8),
	.result_b_8(result_b_8),
	.result_a_7(result_a_7),
	.result_b_7(result_b_7),
	.result_a_6(result_a_6),
	.result_b_6(result_b_6),
	.result_a_5(result_a_5),
	.result_b_5(result_b_5),
	.result_a_4(result_a_4),
	.result_b_4(result_b_4),
	.result_a_3(result_a_3),
	.result_b_3(result_b_3),
	.result_a_2(result_a_2),
	.result_b_2(result_b_2),
	.result_a_1(result_a_1),
	.result_b_1(result_b_1),
	.result_a_0(result_a_0),
	.result_b_0(result_b_0),
	.dffe471(dffe47),
	.dffe241(dffe24),
	.dffe351(dffe35),
	.dffe481(dffe48),
	.dffe251(dffe25),
	.dffe261(dffe26),
	.dffe271(dffe27),
	.dffe281(dffe28),
	.dffe291(dffe29),
	.dffe301(dffe30),
	.dffe311(dffe31),
	.dffe321(dffe32),
	.dffe331(dffe33),
	.dffe341(dffe34),
	.dffe361(dffe36),
	.dffe371(dffe37),
	.dffe381(dffe38),
	.dffe391(dffe39),
	.dffe401(dffe40),
	.dffe411(dffe41),
	.dffe421(dffe42),
	.dffe431(dffe43),
	.dffe441(dffe44),
	.dffe451(dffe45),
	.dffe461(dffe46),
	.clock(clock),
	.clken(clken));

endmodule

module sine_add_sub_5pi (
	result_a_46,
	result_b_46,
	result_a_23,
	result_b_23,
	result_a_34,
	result_b_34,
	result_a_47,
	result_b_47,
	result_a_24,
	result_b_24,
	result_a_25,
	result_b_25,
	result_a_26,
	result_b_26,
	result_a_27,
	result_b_27,
	result_a_28,
	result_b_28,
	result_a_29,
	result_b_29,
	result_a_30,
	result_b_30,
	result_a_31,
	result_b_31,
	result_a_32,
	result_b_32,
	result_a_33,
	result_b_33,
	result_a_35,
	result_b_35,
	result_a_36,
	result_b_36,
	result_a_37,
	result_b_37,
	result_a_38,
	result_b_38,
	result_a_39,
	result_b_39,
	result_a_40,
	result_b_40,
	result_a_41,
	result_b_41,
	result_a_42,
	result_b_42,
	result_a_43,
	result_b_43,
	result_a_44,
	result_b_44,
	result_a_45,
	result_b_45,
	result_a_22,
	result_b_22,
	result_a_21,
	result_b_21,
	result_a_20,
	result_b_20,
	result_a_19,
	result_b_19,
	result_a_18,
	result_b_18,
	result_a_17,
	result_b_17,
	result_a_16,
	result_b_16,
	result_a_15,
	result_b_15,
	result_a_14,
	result_b_14,
	result_a_13,
	result_b_13,
	result_a_12,
	result_b_12,
	result_a_11,
	result_b_11,
	result_a_10,
	result_b_10,
	result_a_9,
	result_b_9,
	result_a_8,
	result_b_8,
	result_a_7,
	result_b_7,
	result_a_6,
	result_b_6,
	result_a_5,
	result_b_5,
	result_a_4,
	result_b_4,
	result_a_3,
	result_b_3,
	result_a_2,
	result_b_2,
	result_a_1,
	result_b_1,
	result_a_0,
	result_b_0,
	dffe471,
	dffe241,
	dffe351,
	dffe481,
	dffe251,
	dffe261,
	dffe271,
	dffe281,
	dffe291,
	dffe301,
	dffe311,
	dffe321,
	dffe331,
	dffe341,
	dffe361,
	dffe371,
	dffe381,
	dffe391,
	dffe401,
	dffe411,
	dffe421,
	dffe431,
	dffe441,
	dffe451,
	dffe461,
	clock,
	clken)/* synthesis synthesis_greybox=1 */;
input 	result_a_46;
input 	result_b_46;
input 	result_a_23;
input 	result_b_23;
input 	result_a_34;
input 	result_b_34;
input 	result_a_47;
input 	result_b_47;
input 	result_a_24;
input 	result_b_24;
input 	result_a_25;
input 	result_b_25;
input 	result_a_26;
input 	result_b_26;
input 	result_a_27;
input 	result_b_27;
input 	result_a_28;
input 	result_b_28;
input 	result_a_29;
input 	result_b_29;
input 	result_a_30;
input 	result_b_30;
input 	result_a_31;
input 	result_b_31;
input 	result_a_32;
input 	result_b_32;
input 	result_a_33;
input 	result_b_33;
input 	result_a_35;
input 	result_b_35;
input 	result_a_36;
input 	result_b_36;
input 	result_a_37;
input 	result_b_37;
input 	result_a_38;
input 	result_b_38;
input 	result_a_39;
input 	result_b_39;
input 	result_a_40;
input 	result_b_40;
input 	result_a_41;
input 	result_b_41;
input 	result_a_42;
input 	result_b_42;
input 	result_a_43;
input 	result_b_43;
input 	result_a_44;
input 	result_b_44;
input 	result_a_45;
input 	result_b_45;
input 	result_a_22;
input 	result_b_22;
input 	result_a_21;
input 	result_b_21;
input 	result_a_20;
input 	result_b_20;
input 	result_a_19;
input 	result_b_19;
input 	result_a_18;
input 	result_b_18;
input 	result_a_17;
input 	result_b_17;
input 	result_a_16;
input 	result_b_16;
input 	result_a_15;
input 	result_b_15;
input 	result_a_14;
input 	result_b_14;
input 	result_a_13;
input 	result_b_13;
input 	result_a_12;
input 	result_b_12;
input 	result_a_11;
input 	result_b_11;
input 	result_a_10;
input 	result_b_10;
input 	result_a_9;
input 	result_b_9;
input 	result_a_8;
input 	result_b_8;
input 	result_a_7;
input 	result_b_7;
input 	result_a_6;
input 	result_b_6;
input 	result_a_5;
input 	result_b_5;
input 	result_a_4;
input 	result_b_4;
input 	result_a_3;
input 	result_b_3;
input 	result_a_2;
input 	result_b_2;
input 	result_a_1;
input 	result_b_1;
input 	result_a_0;
input 	result_b_0;
output 	dffe471;
output 	dffe241;
output 	dffe351;
output 	dffe481;
output 	dffe251;
output 	dffe261;
output 	dffe271;
output 	dffe281;
output 	dffe291;
output 	dffe301;
output 	dffe311;
output 	dffe321;
output 	dffe331;
output 	dffe341;
output 	dffe361;
output 	dffe371;
output 	dffe381;
output 	dffe391;
output 	dffe401;
output 	dffe411;
output 	dffe421;
output 	dffe431;
output 	dffe441;
output 	dffe451;
output 	dffe461;
input 	clock;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~COUT ;
wire \add_sub_cella[18]~COUT ;
wire \add_sub_cella[19]~COUT ;
wire \add_sub_cella[20]~COUT ;
wire \add_sub_cella[21]~COUT ;
wire \add_sub_cella[22]~COUT ;
wire \add_sub_cella[23]~COUT ;
wire \add_sub_cella[24]~COUT ;
wire \add_sub_cella[25]~COUT ;
wire \add_sub_cella[26]~COUT ;
wire \add_sub_cella[27]~COUT ;
wire \add_sub_cella[28]~COUT ;
wire \add_sub_cella[29]~COUT ;
wire \add_sub_cella[30]~COUT ;
wire \add_sub_cella[31]~COUT ;
wire \add_sub_cella[32]~COUT ;
wire \add_sub_cella[33]~COUT ;
wire \add_sub_cella[34]~COUT ;
wire \add_sub_cella[35]~COUT ;
wire \add_sub_cella[36]~COUT ;
wire \add_sub_cella[37]~COUT ;
wire \add_sub_cella[38]~COUT ;
wire \add_sub_cella[39]~COUT ;
wire \add_sub_cella[40]~COUT ;
wire \add_sub_cella[41]~COUT ;
wire \add_sub_cella[42]~COUT ;
wire \add_sub_cella[43]~COUT ;
wire \add_sub_cella[44]~COUT ;
wire \add_sub_cella[45]~COUT ;
wire \add_sub_cella[46]~sumout ;
wire \add_sub_cella[23]~sumout ;
wire \add_sub_cella[34]~sumout ;
wire \add_sub_cella[46]~COUT ;
wire \add_sub_cella[47]~sumout ;
wire \add_sub_cella[24]~sumout ;
wire \add_sub_cella[25]~sumout ;
wire \add_sub_cella[26]~sumout ;
wire \add_sub_cella[27]~sumout ;
wire \add_sub_cella[28]~sumout ;
wire \add_sub_cella[29]~sumout ;
wire \add_sub_cella[30]~sumout ;
wire \add_sub_cella[31]~sumout ;
wire \add_sub_cella[32]~sumout ;
wire \add_sub_cella[33]~sumout ;
wire \add_sub_cella[35]~sumout ;
wire \add_sub_cella[36]~sumout ;
wire \add_sub_cella[37]~sumout ;
wire \add_sub_cella[38]~sumout ;
wire \add_sub_cella[39]~sumout ;
wire \add_sub_cella[40]~sumout ;
wire \add_sub_cella[41]~sumout ;
wire \add_sub_cella[42]~sumout ;
wire \add_sub_cella[43]~sumout ;
wire \add_sub_cella[44]~sumout ;
wire \add_sub_cella[45]~sumout ;


dffeas dffe47(
	.clk(clock),
	.d(\add_sub_cella[46]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe471),
	.prn(vcc));
defparam dffe47.is_wysiwyg = "true";
defparam dffe47.power_up = "low";

dffeas dffe24(
	.clk(clock),
	.d(\add_sub_cella[23]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe241),
	.prn(vcc));
defparam dffe24.is_wysiwyg = "true";
defparam dffe24.power_up = "low";

dffeas dffe35(
	.clk(clock),
	.d(\add_sub_cella[34]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe351),
	.prn(vcc));
defparam dffe35.is_wysiwyg = "true";
defparam dffe35.power_up = "low";

dffeas dffe48(
	.clk(clock),
	.d(\add_sub_cella[47]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe481),
	.prn(vcc));
defparam dffe48.is_wysiwyg = "true";
defparam dffe48.power_up = "low";

dffeas dffe25(
	.clk(clock),
	.d(\add_sub_cella[24]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe251),
	.prn(vcc));
defparam dffe25.is_wysiwyg = "true";
defparam dffe25.power_up = "low";

dffeas dffe26(
	.clk(clock),
	.d(\add_sub_cella[25]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe261),
	.prn(vcc));
defparam dffe26.is_wysiwyg = "true";
defparam dffe26.power_up = "low";

dffeas dffe27(
	.clk(clock),
	.d(\add_sub_cella[26]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe271),
	.prn(vcc));
defparam dffe27.is_wysiwyg = "true";
defparam dffe27.power_up = "low";

dffeas dffe28(
	.clk(clock),
	.d(\add_sub_cella[27]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe281),
	.prn(vcc));
defparam dffe28.is_wysiwyg = "true";
defparam dffe28.power_up = "low";

dffeas dffe29(
	.clk(clock),
	.d(\add_sub_cella[28]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe291),
	.prn(vcc));
defparam dffe29.is_wysiwyg = "true";
defparam dffe29.power_up = "low";

dffeas dffe30(
	.clk(clock),
	.d(\add_sub_cella[29]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe301),
	.prn(vcc));
defparam dffe30.is_wysiwyg = "true";
defparam dffe30.power_up = "low";

dffeas dffe31(
	.clk(clock),
	.d(\add_sub_cella[30]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe311),
	.prn(vcc));
defparam dffe31.is_wysiwyg = "true";
defparam dffe31.power_up = "low";

dffeas dffe32(
	.clk(clock),
	.d(\add_sub_cella[31]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe321),
	.prn(vcc));
defparam dffe32.is_wysiwyg = "true";
defparam dffe32.power_up = "low";

dffeas dffe33(
	.clk(clock),
	.d(\add_sub_cella[32]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe331),
	.prn(vcc));
defparam dffe33.is_wysiwyg = "true";
defparam dffe33.power_up = "low";

dffeas dffe34(
	.clk(clock),
	.d(\add_sub_cella[33]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe341),
	.prn(vcc));
defparam dffe34.is_wysiwyg = "true";
defparam dffe34.power_up = "low";

dffeas dffe36(
	.clk(clock),
	.d(\add_sub_cella[35]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe361),
	.prn(vcc));
defparam dffe36.is_wysiwyg = "true";
defparam dffe36.power_up = "low";

dffeas dffe37(
	.clk(clock),
	.d(\add_sub_cella[36]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe371),
	.prn(vcc));
defparam dffe37.is_wysiwyg = "true";
defparam dffe37.power_up = "low";

dffeas dffe38(
	.clk(clock),
	.d(\add_sub_cella[37]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe381),
	.prn(vcc));
defparam dffe38.is_wysiwyg = "true";
defparam dffe38.power_up = "low";

dffeas dffe39(
	.clk(clock),
	.d(\add_sub_cella[38]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe391),
	.prn(vcc));
defparam dffe39.is_wysiwyg = "true";
defparam dffe39.power_up = "low";

dffeas dffe40(
	.clk(clock),
	.d(\add_sub_cella[39]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe401),
	.prn(vcc));
defparam dffe40.is_wysiwyg = "true";
defparam dffe40.power_up = "low";

dffeas dffe41(
	.clk(clock),
	.d(\add_sub_cella[40]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe411),
	.prn(vcc));
defparam dffe41.is_wysiwyg = "true";
defparam dffe41.power_up = "low";

dffeas dffe42(
	.clk(clock),
	.d(\add_sub_cella[41]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe421),
	.prn(vcc));
defparam dffe42.is_wysiwyg = "true";
defparam dffe42.power_up = "low";

dffeas dffe43(
	.clk(clock),
	.d(\add_sub_cella[42]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe431),
	.prn(vcc));
defparam dffe43.is_wysiwyg = "true";
defparam dffe43.power_up = "low";

dffeas dffe44(
	.clk(clock),
	.d(\add_sub_cella[43]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe441),
	.prn(vcc));
defparam dffe44.is_wysiwyg = "true";
defparam dffe44.power_up = "low";

dffeas dffe45(
	.clk(clock),
	.d(\add_sub_cella[44]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe451),
	.prn(vcc));
defparam dffe45.is_wysiwyg = "true";
defparam dffe45.power_up = "low";

dffeas dffe46(
	.clk(clock),
	.d(\add_sub_cella[45]~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe461),
	.prn(vcc));
defparam dffe46.is_wysiwyg = "true";
defparam dffe46.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_0),
	.datae(gnd),
	.dataf(!result_b_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_1),
	.datae(gnd),
	.dataf(!result_b_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_2),
	.datae(gnd),
	.dataf(!result_b_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_3),
	.datae(gnd),
	.dataf(!result_b_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_4),
	.datae(gnd),
	.dataf(!result_b_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_5),
	.datae(gnd),
	.dataf(!result_b_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_6),
	.datae(gnd),
	.dataf(!result_b_6),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_7),
	.datae(gnd),
	.dataf(!result_b_7),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_8),
	.datae(gnd),
	.dataf(!result_b_8),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_9),
	.datae(gnd),
	.dataf(!result_b_9),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_10),
	.datae(gnd),
	.dataf(!result_b_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_11),
	.datae(gnd),
	.dataf(!result_b_11),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_12),
	.datae(gnd),
	.dataf(!result_b_12),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_13),
	.datae(gnd),
	.dataf(!result_b_13),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_14),
	.datae(gnd),
	.dataf(!result_b_14),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_15),
	.datae(gnd),
	.dataf(!result_b_15),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_16),
	.datae(gnd),
	.dataf(!result_b_16),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_17),
	.datae(gnd),
	.dataf(!result_b_17),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[17]~COUT ),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[18] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_18),
	.datae(gnd),
	.dataf(!result_b_18),
	.datag(gnd),
	.cin(\add_sub_cella[17]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[18]~COUT ),
	.shareout());
defparam \add_sub_cella[18] .extended_lut = "off";
defparam \add_sub_cella[18] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[18] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[19] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_19),
	.datae(gnd),
	.dataf(!result_b_19),
	.datag(gnd),
	.cin(\add_sub_cella[18]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[19]~COUT ),
	.shareout());
defparam \add_sub_cella[19] .extended_lut = "off";
defparam \add_sub_cella[19] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[19] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[20] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_20),
	.datae(gnd),
	.dataf(!result_b_20),
	.datag(gnd),
	.cin(\add_sub_cella[19]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[20]~COUT ),
	.shareout());
defparam \add_sub_cella[20] .extended_lut = "off";
defparam \add_sub_cella[20] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[20] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[21] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_21),
	.datae(gnd),
	.dataf(!result_b_21),
	.datag(gnd),
	.cin(\add_sub_cella[20]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[21]~COUT ),
	.shareout());
defparam \add_sub_cella[21] .extended_lut = "off";
defparam \add_sub_cella[21] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[21] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[22] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_22),
	.datae(gnd),
	.dataf(!result_b_22),
	.datag(gnd),
	.cin(\add_sub_cella[21]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[22]~COUT ),
	.shareout());
defparam \add_sub_cella[22] .extended_lut = "off";
defparam \add_sub_cella[22] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[22] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[23] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_23),
	.datae(gnd),
	.dataf(!result_b_23),
	.datag(gnd),
	.cin(\add_sub_cella[22]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[23]~sumout ),
	.cout(\add_sub_cella[23]~COUT ),
	.shareout());
defparam \add_sub_cella[23] .extended_lut = "off";
defparam \add_sub_cella[23] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[23] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[24] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_24),
	.datae(gnd),
	.dataf(!result_b_24),
	.datag(gnd),
	.cin(\add_sub_cella[23]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[24]~sumout ),
	.cout(\add_sub_cella[24]~COUT ),
	.shareout());
defparam \add_sub_cella[24] .extended_lut = "off";
defparam \add_sub_cella[24] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[24] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[25] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_25),
	.datae(gnd),
	.dataf(!result_b_25),
	.datag(gnd),
	.cin(\add_sub_cella[24]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[25]~sumout ),
	.cout(\add_sub_cella[25]~COUT ),
	.shareout());
defparam \add_sub_cella[25] .extended_lut = "off";
defparam \add_sub_cella[25] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[25] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[26] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_26),
	.datae(gnd),
	.dataf(!result_b_26),
	.datag(gnd),
	.cin(\add_sub_cella[25]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[26]~sumout ),
	.cout(\add_sub_cella[26]~COUT ),
	.shareout());
defparam \add_sub_cella[26] .extended_lut = "off";
defparam \add_sub_cella[26] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[26] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[27] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_27),
	.datae(gnd),
	.dataf(!result_b_27),
	.datag(gnd),
	.cin(\add_sub_cella[26]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[27]~sumout ),
	.cout(\add_sub_cella[27]~COUT ),
	.shareout());
defparam \add_sub_cella[27] .extended_lut = "off";
defparam \add_sub_cella[27] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[27] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[28] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_28),
	.datae(gnd),
	.dataf(!result_b_28),
	.datag(gnd),
	.cin(\add_sub_cella[27]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[28]~sumout ),
	.cout(\add_sub_cella[28]~COUT ),
	.shareout());
defparam \add_sub_cella[28] .extended_lut = "off";
defparam \add_sub_cella[28] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[28] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[29] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_29),
	.datae(gnd),
	.dataf(!result_b_29),
	.datag(gnd),
	.cin(\add_sub_cella[28]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[29]~sumout ),
	.cout(\add_sub_cella[29]~COUT ),
	.shareout());
defparam \add_sub_cella[29] .extended_lut = "off";
defparam \add_sub_cella[29] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[29] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[30] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_30),
	.datae(gnd),
	.dataf(!result_b_30),
	.datag(gnd),
	.cin(\add_sub_cella[29]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[30]~sumout ),
	.cout(\add_sub_cella[30]~COUT ),
	.shareout());
defparam \add_sub_cella[30] .extended_lut = "off";
defparam \add_sub_cella[30] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[30] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[31] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_31),
	.datae(gnd),
	.dataf(!result_b_31),
	.datag(gnd),
	.cin(\add_sub_cella[30]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[31]~sumout ),
	.cout(\add_sub_cella[31]~COUT ),
	.shareout());
defparam \add_sub_cella[31] .extended_lut = "off";
defparam \add_sub_cella[31] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[31] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[32] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_32),
	.datae(gnd),
	.dataf(!result_b_32),
	.datag(gnd),
	.cin(\add_sub_cella[31]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[32]~sumout ),
	.cout(\add_sub_cella[32]~COUT ),
	.shareout());
defparam \add_sub_cella[32] .extended_lut = "off";
defparam \add_sub_cella[32] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[32] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[33] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_33),
	.datae(gnd),
	.dataf(!result_b_33),
	.datag(gnd),
	.cin(\add_sub_cella[32]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[33]~sumout ),
	.cout(\add_sub_cella[33]~COUT ),
	.shareout());
defparam \add_sub_cella[33] .extended_lut = "off";
defparam \add_sub_cella[33] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[33] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[34] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_34),
	.datae(gnd),
	.dataf(!result_b_34),
	.datag(gnd),
	.cin(\add_sub_cella[33]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[34]~sumout ),
	.cout(\add_sub_cella[34]~COUT ),
	.shareout());
defparam \add_sub_cella[34] .extended_lut = "off";
defparam \add_sub_cella[34] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[34] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[35] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_35),
	.datae(gnd),
	.dataf(!result_b_35),
	.datag(gnd),
	.cin(\add_sub_cella[34]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[35]~sumout ),
	.cout(\add_sub_cella[35]~COUT ),
	.shareout());
defparam \add_sub_cella[35] .extended_lut = "off";
defparam \add_sub_cella[35] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[35] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[36] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_36),
	.datae(gnd),
	.dataf(!result_b_36),
	.datag(gnd),
	.cin(\add_sub_cella[35]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[36]~sumout ),
	.cout(\add_sub_cella[36]~COUT ),
	.shareout());
defparam \add_sub_cella[36] .extended_lut = "off";
defparam \add_sub_cella[36] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[36] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[37] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_37),
	.datae(gnd),
	.dataf(!result_b_37),
	.datag(gnd),
	.cin(\add_sub_cella[36]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[37]~sumout ),
	.cout(\add_sub_cella[37]~COUT ),
	.shareout());
defparam \add_sub_cella[37] .extended_lut = "off";
defparam \add_sub_cella[37] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[37] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[38] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_38),
	.datae(gnd),
	.dataf(!result_b_38),
	.datag(gnd),
	.cin(\add_sub_cella[37]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[38]~sumout ),
	.cout(\add_sub_cella[38]~COUT ),
	.shareout());
defparam \add_sub_cella[38] .extended_lut = "off";
defparam \add_sub_cella[38] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[38] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[39] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_39),
	.datae(gnd),
	.dataf(!result_b_39),
	.datag(gnd),
	.cin(\add_sub_cella[38]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[39]~sumout ),
	.cout(\add_sub_cella[39]~COUT ),
	.shareout());
defparam \add_sub_cella[39] .extended_lut = "off";
defparam \add_sub_cella[39] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[39] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[40] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_40),
	.datae(gnd),
	.dataf(!result_b_40),
	.datag(gnd),
	.cin(\add_sub_cella[39]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[40]~sumout ),
	.cout(\add_sub_cella[40]~COUT ),
	.shareout());
defparam \add_sub_cella[40] .extended_lut = "off";
defparam \add_sub_cella[40] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[40] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[41] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_41),
	.datae(gnd),
	.dataf(!result_b_41),
	.datag(gnd),
	.cin(\add_sub_cella[40]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[41]~sumout ),
	.cout(\add_sub_cella[41]~COUT ),
	.shareout());
defparam \add_sub_cella[41] .extended_lut = "off";
defparam \add_sub_cella[41] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[41] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[42] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_42),
	.datae(gnd),
	.dataf(!result_b_42),
	.datag(gnd),
	.cin(\add_sub_cella[41]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[42]~sumout ),
	.cout(\add_sub_cella[42]~COUT ),
	.shareout());
defparam \add_sub_cella[42] .extended_lut = "off";
defparam \add_sub_cella[42] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[42] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[43] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_43),
	.datae(gnd),
	.dataf(!result_b_43),
	.datag(gnd),
	.cin(\add_sub_cella[42]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[43]~sumout ),
	.cout(\add_sub_cella[43]~COUT ),
	.shareout());
defparam \add_sub_cella[43] .extended_lut = "off";
defparam \add_sub_cella[43] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[43] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[44] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_44),
	.datae(gnd),
	.dataf(!result_b_44),
	.datag(gnd),
	.cin(\add_sub_cella[43]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[44]~sumout ),
	.cout(\add_sub_cella[44]~COUT ),
	.shareout());
defparam \add_sub_cella[44] .extended_lut = "off";
defparam \add_sub_cella[44] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[44] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[45] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_45),
	.datae(gnd),
	.dataf(!result_b_45),
	.datag(gnd),
	.cin(\add_sub_cella[44]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[45]~sumout ),
	.cout(\add_sub_cella[45]~COUT ),
	.shareout());
defparam \add_sub_cella[45] .extended_lut = "off";
defparam \add_sub_cella[45] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[45] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[46] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_46),
	.datae(gnd),
	.dataf(!result_b_46),
	.datag(gnd),
	.cin(\add_sub_cella[45]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[46]~sumout ),
	.cout(\add_sub_cella[46]~COUT ),
	.shareout());
defparam \add_sub_cella[46] .extended_lut = "off";
defparam \add_sub_cella[46] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[46] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[47] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_a_47),
	.datae(gnd),
	.dataf(!result_b_47),
	.datag(gnd),
	.cin(\add_sub_cella[46]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[47]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[47] .extended_lut = "off";
defparam \add_sub_cella[47] .lut_mask = 64'h0000FF00000000FF;
defparam \add_sub_cella[47] .shared_arith = "off";

endmodule

module sine_lmsd (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	q_a_10,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	q_a_16,
	q_a_17,
	q_a_18,
	q_a_19,
	q_a_20,
	q_a_21,
	q_a_22,
	q_a_23,
	q_a_01,
	q_a_110,
	q_a_24,
	q_a_31,
	q_a_41,
	q_a_51,
	q_a_61,
	q_a_71,
	q_a_81,
	q_a_91,
	q_a_101,
	q_a_111,
	q_a_121,
	q_a_131,
	q_a_141,
	q_a_151,
	q_a_161,
	q_a_171,
	q_a_181,
	q_a_191,
	q_a_201,
	q_a_211,
	q_a_221,
	q_a_231,
	result_output_reg_46,
	result_output_reg_23,
	result_output_reg_34,
	result_output_reg_47,
	result_output_reg_24,
	result_output_reg_25,
	result_output_reg_26,
	result_output_reg_27,
	result_output_reg_28,
	result_output_reg_29,
	result_output_reg_30,
	result_output_reg_31,
	result_output_reg_32,
	result_output_reg_33,
	result_output_reg_35,
	result_output_reg_36,
	result_output_reg_37,
	result_output_reg_38,
	result_output_reg_39,
	result_output_reg_40,
	result_output_reg_41,
	result_output_reg_42,
	result_output_reg_43,
	result_output_reg_44,
	result_output_reg_45,
	result_output_reg_22,
	result_output_reg_21,
	result_output_reg_20,
	result_output_reg_19,
	result_output_reg_18,
	result_output_reg_17,
	result_output_reg_16,
	result_output_reg_15,
	result_output_reg_14,
	result_output_reg_13,
	result_output_reg_12,
	result_output_reg_11,
	result_output_reg_10,
	result_output_reg_9,
	result_output_reg_8,
	result_output_reg_7,
	result_output_reg_6,
	result_output_reg_5,
	result_output_reg_4,
	result_output_reg_3,
	result_output_reg_2,
	result_output_reg_1,
	result_output_reg_0,
	clk,
	clken)/* synthesis synthesis_greybox=1 */;
input 	q_a_0;
input 	q_a_1;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_5;
input 	q_a_6;
input 	q_a_7;
input 	q_a_8;
input 	q_a_9;
input 	q_a_10;
input 	q_a_11;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_15;
input 	q_a_16;
input 	q_a_17;
input 	q_a_18;
input 	q_a_19;
input 	q_a_20;
input 	q_a_21;
input 	q_a_22;
input 	q_a_23;
input 	q_a_01;
input 	q_a_110;
input 	q_a_24;
input 	q_a_31;
input 	q_a_41;
input 	q_a_51;
input 	q_a_61;
input 	q_a_71;
input 	q_a_81;
input 	q_a_91;
input 	q_a_101;
input 	q_a_111;
input 	q_a_121;
input 	q_a_131;
input 	q_a_141;
input 	q_a_151;
input 	q_a_161;
input 	q_a_171;
input 	q_a_181;
input 	q_a_191;
input 	q_a_201;
input 	q_a_211;
input 	q_a_221;
input 	q_a_231;
output 	result_output_reg_46;
output 	result_output_reg_23;
output 	result_output_reg_34;
output 	result_output_reg_47;
output 	result_output_reg_24;
output 	result_output_reg_25;
output 	result_output_reg_26;
output 	result_output_reg_27;
output 	result_output_reg_28;
output 	result_output_reg_29;
output 	result_output_reg_30;
output 	result_output_reg_31;
output 	result_output_reg_32;
output 	result_output_reg_33;
output 	result_output_reg_35;
output 	result_output_reg_36;
output 	result_output_reg_37;
output 	result_output_reg_38;
output 	result_output_reg_39;
output 	result_output_reg_40;
output 	result_output_reg_41;
output 	result_output_reg_42;
output 	result_output_reg_43;
output 	result_output_reg_44;
output 	result_output_reg_45;
output 	result_output_reg_22;
output 	result_output_reg_21;
output 	result_output_reg_20;
output 	result_output_reg_19;
output 	result_output_reg_18;
output 	result_output_reg_17;
output 	result_output_reg_16;
output 	result_output_reg_15;
output 	result_output_reg_14;
output 	result_output_reg_13;
output 	result_output_reg_12;
output 	result_output_reg_11;
output 	result_output_reg_10;
output 	result_output_reg_9;
output 	result_output_reg_8;
output 	result_output_reg_7;
output 	result_output_reg_6;
output 	result_output_reg_5;
output 	result_output_reg_4;
output 	result_output_reg_3;
output 	result_output_reg_2;
output 	result_output_reg_1;
output 	result_output_reg_0;
input 	clk;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_lpm_mult_1 lpm_mult_component(
	.dataa({q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.datab({q_a_231,q_a_221,q_a_211,q_a_201,q_a_191,q_a_181,q_a_171,q_a_161,q_a_151,q_a_141,q_a_131,q_a_121,q_a_111,q_a_101,q_a_91,q_a_81,q_a_71,q_a_61,q_a_51,q_a_41,q_a_31,q_a_24,q_a_110,q_a_01}),
	.result_output_reg_46(result_output_reg_46),
	.result_output_reg_23(result_output_reg_23),
	.result_output_reg_34(result_output_reg_34),
	.result_output_reg_47(result_output_reg_47),
	.result_output_reg_24(result_output_reg_24),
	.result_output_reg_25(result_output_reg_25),
	.result_output_reg_26(result_output_reg_26),
	.result_output_reg_27(result_output_reg_27),
	.result_output_reg_28(result_output_reg_28),
	.result_output_reg_29(result_output_reg_29),
	.result_output_reg_30(result_output_reg_30),
	.result_output_reg_31(result_output_reg_31),
	.result_output_reg_32(result_output_reg_32),
	.result_output_reg_33(result_output_reg_33),
	.result_output_reg_35(result_output_reg_35),
	.result_output_reg_36(result_output_reg_36),
	.result_output_reg_37(result_output_reg_37),
	.result_output_reg_38(result_output_reg_38),
	.result_output_reg_39(result_output_reg_39),
	.result_output_reg_40(result_output_reg_40),
	.result_output_reg_41(result_output_reg_41),
	.result_output_reg_42(result_output_reg_42),
	.result_output_reg_43(result_output_reg_43),
	.result_output_reg_44(result_output_reg_44),
	.result_output_reg_45(result_output_reg_45),
	.result_output_reg_22(result_output_reg_22),
	.result_output_reg_21(result_output_reg_21),
	.result_output_reg_20(result_output_reg_20),
	.result_output_reg_19(result_output_reg_19),
	.result_output_reg_18(result_output_reg_18),
	.result_output_reg_17(result_output_reg_17),
	.result_output_reg_16(result_output_reg_16),
	.result_output_reg_15(result_output_reg_15),
	.result_output_reg_14(result_output_reg_14),
	.result_output_reg_13(result_output_reg_13),
	.result_output_reg_12(result_output_reg_12),
	.result_output_reg_11(result_output_reg_11),
	.result_output_reg_10(result_output_reg_10),
	.result_output_reg_9(result_output_reg_9),
	.result_output_reg_8(result_output_reg_8),
	.result_output_reg_7(result_output_reg_7),
	.result_output_reg_6(result_output_reg_6),
	.result_output_reg_5(result_output_reg_5),
	.result_output_reg_4(result_output_reg_4),
	.result_output_reg_3(result_output_reg_3),
	.result_output_reg_2(result_output_reg_2),
	.result_output_reg_1(result_output_reg_1),
	.result_output_reg_0(result_output_reg_0),
	.clock(clk),
	.clken(clken));

endmodule

module sine_lpm_mult_1 (
	dataa,
	datab,
	result_output_reg_46,
	result_output_reg_23,
	result_output_reg_34,
	result_output_reg_47,
	result_output_reg_24,
	result_output_reg_25,
	result_output_reg_26,
	result_output_reg_27,
	result_output_reg_28,
	result_output_reg_29,
	result_output_reg_30,
	result_output_reg_31,
	result_output_reg_32,
	result_output_reg_33,
	result_output_reg_35,
	result_output_reg_36,
	result_output_reg_37,
	result_output_reg_38,
	result_output_reg_39,
	result_output_reg_40,
	result_output_reg_41,
	result_output_reg_42,
	result_output_reg_43,
	result_output_reg_44,
	result_output_reg_45,
	result_output_reg_22,
	result_output_reg_21,
	result_output_reg_20,
	result_output_reg_19,
	result_output_reg_18,
	result_output_reg_17,
	result_output_reg_16,
	result_output_reg_15,
	result_output_reg_14,
	result_output_reg_13,
	result_output_reg_12,
	result_output_reg_11,
	result_output_reg_10,
	result_output_reg_9,
	result_output_reg_8,
	result_output_reg_7,
	result_output_reg_6,
	result_output_reg_5,
	result_output_reg_4,
	result_output_reg_3,
	result_output_reg_2,
	result_output_reg_1,
	result_output_reg_0,
	clock,
	clken)/* synthesis synthesis_greybox=1 */;
input 	[23:0] dataa;
input 	[23:0] datab;
output 	result_output_reg_46;
output 	result_output_reg_23;
output 	result_output_reg_34;
output 	result_output_reg_47;
output 	result_output_reg_24;
output 	result_output_reg_25;
output 	result_output_reg_26;
output 	result_output_reg_27;
output 	result_output_reg_28;
output 	result_output_reg_29;
output 	result_output_reg_30;
output 	result_output_reg_31;
output 	result_output_reg_32;
output 	result_output_reg_33;
output 	result_output_reg_35;
output 	result_output_reg_36;
output 	result_output_reg_37;
output 	result_output_reg_38;
output 	result_output_reg_39;
output 	result_output_reg_40;
output 	result_output_reg_41;
output 	result_output_reg_42;
output 	result_output_reg_43;
output 	result_output_reg_44;
output 	result_output_reg_45;
output 	result_output_reg_22;
output 	result_output_reg_21;
output 	result_output_reg_20;
output 	result_output_reg_19;
output 	result_output_reg_18;
output 	result_output_reg_17;
output 	result_output_reg_16;
output 	result_output_reg_15;
output 	result_output_reg_14;
output 	result_output_reg_13;
output 	result_output_reg_12;
output 	result_output_reg_11;
output 	result_output_reg_10;
output 	result_output_reg_9;
output 	result_output_reg_8;
output 	result_output_reg_7;
output 	result_output_reg_6;
output 	result_output_reg_5;
output 	result_output_reg_4;
output 	result_output_reg_3;
output 	result_output_reg_2;
output 	result_output_reg_1;
output 	result_output_reg_0;
input 	clock;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_mult_5cu auto_generated(
	.dataa({dataa[23],dataa[22],dataa[21],dataa[20],dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({datab[23],datab[22],datab[21],datab[20],datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.result_output_reg_46(result_output_reg_46),
	.result_output_reg_23(result_output_reg_23),
	.result_output_reg_34(result_output_reg_34),
	.result_output_reg_47(result_output_reg_47),
	.result_output_reg_24(result_output_reg_24),
	.result_output_reg_25(result_output_reg_25),
	.result_output_reg_26(result_output_reg_26),
	.result_output_reg_27(result_output_reg_27),
	.result_output_reg_28(result_output_reg_28),
	.result_output_reg_29(result_output_reg_29),
	.result_output_reg_30(result_output_reg_30),
	.result_output_reg_31(result_output_reg_31),
	.result_output_reg_32(result_output_reg_32),
	.result_output_reg_33(result_output_reg_33),
	.result_output_reg_35(result_output_reg_35),
	.result_output_reg_36(result_output_reg_36),
	.result_output_reg_37(result_output_reg_37),
	.result_output_reg_38(result_output_reg_38),
	.result_output_reg_39(result_output_reg_39),
	.result_output_reg_40(result_output_reg_40),
	.result_output_reg_41(result_output_reg_41),
	.result_output_reg_42(result_output_reg_42),
	.result_output_reg_43(result_output_reg_43),
	.result_output_reg_44(result_output_reg_44),
	.result_output_reg_45(result_output_reg_45),
	.result_output_reg_22(result_output_reg_22),
	.result_output_reg_21(result_output_reg_21),
	.result_output_reg_20(result_output_reg_20),
	.result_output_reg_19(result_output_reg_19),
	.result_output_reg_18(result_output_reg_18),
	.result_output_reg_17(result_output_reg_17),
	.result_output_reg_16(result_output_reg_16),
	.result_output_reg_15(result_output_reg_15),
	.result_output_reg_14(result_output_reg_14),
	.result_output_reg_13(result_output_reg_13),
	.result_output_reg_12(result_output_reg_12),
	.result_output_reg_11(result_output_reg_11),
	.result_output_reg_10(result_output_reg_10),
	.result_output_reg_9(result_output_reg_9),
	.result_output_reg_8(result_output_reg_8),
	.result_output_reg_7(result_output_reg_7),
	.result_output_reg_6(result_output_reg_6),
	.result_output_reg_5(result_output_reg_5),
	.result_output_reg_4(result_output_reg_4),
	.result_output_reg_3(result_output_reg_3),
	.result_output_reg_2(result_output_reg_2),
	.result_output_reg_1(result_output_reg_1),
	.result_output_reg_0(result_output_reg_0),
	.clock(clock),
	.clken(clken));

endmodule

module sine_mult_5cu (
	dataa,
	datab,
	result_output_reg_46,
	result_output_reg_23,
	result_output_reg_34,
	result_output_reg_47,
	result_output_reg_24,
	result_output_reg_25,
	result_output_reg_26,
	result_output_reg_27,
	result_output_reg_28,
	result_output_reg_29,
	result_output_reg_30,
	result_output_reg_31,
	result_output_reg_32,
	result_output_reg_33,
	result_output_reg_35,
	result_output_reg_36,
	result_output_reg_37,
	result_output_reg_38,
	result_output_reg_39,
	result_output_reg_40,
	result_output_reg_41,
	result_output_reg_42,
	result_output_reg_43,
	result_output_reg_44,
	result_output_reg_45,
	result_output_reg_22,
	result_output_reg_21,
	result_output_reg_20,
	result_output_reg_19,
	result_output_reg_18,
	result_output_reg_17,
	result_output_reg_16,
	result_output_reg_15,
	result_output_reg_14,
	result_output_reg_13,
	result_output_reg_12,
	result_output_reg_11,
	result_output_reg_10,
	result_output_reg_9,
	result_output_reg_8,
	result_output_reg_7,
	result_output_reg_6,
	result_output_reg_5,
	result_output_reg_4,
	result_output_reg_3,
	result_output_reg_2,
	result_output_reg_1,
	result_output_reg_0,
	clock,
	clken)/* synthesis synthesis_greybox=1 */;
input 	[23:0] dataa;
input 	[23:0] datab;
output 	result_output_reg_46;
output 	result_output_reg_23;
output 	result_output_reg_34;
output 	result_output_reg_47;
output 	result_output_reg_24;
output 	result_output_reg_25;
output 	result_output_reg_26;
output 	result_output_reg_27;
output 	result_output_reg_28;
output 	result_output_reg_29;
output 	result_output_reg_30;
output 	result_output_reg_31;
output 	result_output_reg_32;
output 	result_output_reg_33;
output 	result_output_reg_35;
output 	result_output_reg_36;
output 	result_output_reg_37;
output 	result_output_reg_38;
output 	result_output_reg_39;
output 	result_output_reg_40;
output 	result_output_reg_41;
output 	result_output_reg_42;
output 	result_output_reg_43;
output 	result_output_reg_44;
output 	result_output_reg_45;
output 	result_output_reg_22;
output 	result_output_reg_21;
output 	result_output_reg_20;
output 	result_output_reg_19;
output 	result_output_reg_18;
output 	result_output_reg_17;
output 	result_output_reg_16;
output 	result_output_reg_15;
output 	result_output_reg_14;
output 	result_output_reg_13;
output 	result_output_reg_12;
output 	result_output_reg_11;
output 	result_output_reg_10;
output 	result_output_reg_9;
output 	result_output_reg_8;
output 	result_output_reg_7;
output 	result_output_reg_6;
output 	result_output_reg_5;
output 	result_output_reg_4;
output 	result_output_reg_3;
output 	result_output_reg_2;
output 	result_output_reg_1;
output 	result_output_reg_0;
input 	clock;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mult0~8 ;
wire \Mult0~9 ;
wire \Mult0~10 ;
wire \Mult0~11 ;
wire \Mult0~12 ;
wire \Mult0~13 ;
wire \Mult0~14 ;
wire \Mult0~15 ;
wire \Mult0~16 ;
wire \Mult0~17 ;
wire \Mult0~18 ;
wire \Mult0~19 ;
wire \Mult0~20 ;
wire \Mult0~21 ;
wire \Mult0~22 ;
wire \Mult0~23 ;
wire \dataa_input_reg[0]~q ;
wire \dataa_input_reg[1]~q ;
wire \dataa_input_reg[2]~q ;
wire \dataa_input_reg[3]~q ;
wire \dataa_input_reg[4]~q ;
wire \dataa_input_reg[5]~q ;
wire \dataa_input_reg[6]~q ;
wire \dataa_input_reg[7]~q ;
wire \dataa_input_reg[8]~q ;
wire \dataa_input_reg[9]~q ;
wire \dataa_input_reg[10]~q ;
wire \dataa_input_reg[11]~q ;
wire \dataa_input_reg[12]~q ;
wire \dataa_input_reg[13]~q ;
wire \dataa_input_reg[14]~q ;
wire \dataa_input_reg[15]~q ;
wire \dataa_input_reg[16]~q ;
wire \dataa_input_reg[17]~q ;
wire \dataa_input_reg[18]~q ;
wire \dataa_input_reg[19]~q ;
wire \dataa_input_reg[20]~q ;
wire \dataa_input_reg[21]~q ;
wire \dataa_input_reg[22]~q ;
wire \dataa_input_reg[23]~q ;
wire \datab_input_reg[0]~q ;
wire \datab_input_reg[1]~q ;
wire \datab_input_reg[2]~q ;
wire \datab_input_reg[3]~q ;
wire \datab_input_reg[4]~q ;
wire \datab_input_reg[5]~q ;
wire \datab_input_reg[6]~q ;
wire \datab_input_reg[7]~q ;
wire \datab_input_reg[8]~q ;
wire \datab_input_reg[9]~q ;
wire \datab_input_reg[10]~q ;
wire \datab_input_reg[11]~q ;
wire \datab_input_reg[12]~q ;
wire \datab_input_reg[13]~q ;
wire \datab_input_reg[14]~q ;
wire \datab_input_reg[15]~q ;
wire \datab_input_reg[16]~q ;
wire \datab_input_reg[17]~q ;
wire \datab_input_reg[18]~q ;
wire \datab_input_reg[19]~q ;
wire \datab_input_reg[20]~q ;
wire \datab_input_reg[21]~q ;
wire \datab_input_reg[22]~q ;
wire \datab_input_reg[23]~q ;
wire \result_wire[46] ;
wire \result_extra0_reg[46]~q ;
wire \result_wire[23] ;
wire \result_extra0_reg[23]~q ;
wire \result_wire[34] ;
wire \result_extra0_reg[34]~q ;
wire \result_wire[47] ;
wire \result_extra0_reg[47]~q ;
wire \result_wire[24] ;
wire \result_extra0_reg[24]~q ;
wire \result_wire[25] ;
wire \result_extra0_reg[25]~q ;
wire \result_wire[26] ;
wire \result_extra0_reg[26]~q ;
wire \result_wire[27] ;
wire \result_extra0_reg[27]~q ;
wire \result_wire[28] ;
wire \result_extra0_reg[28]~q ;
wire \result_wire[29] ;
wire \result_extra0_reg[29]~q ;
wire \result_wire[30] ;
wire \result_extra0_reg[30]~q ;
wire \result_wire[31] ;
wire \result_extra0_reg[31]~q ;
wire \result_wire[32] ;
wire \result_extra0_reg[32]~q ;
wire \result_wire[33] ;
wire \result_extra0_reg[33]~q ;
wire \result_wire[35] ;
wire \result_extra0_reg[35]~q ;
wire \result_wire[36] ;
wire \result_extra0_reg[36]~q ;
wire \result_wire[37] ;
wire \result_extra0_reg[37]~q ;
wire \result_wire[38] ;
wire \result_extra0_reg[38]~q ;
wire \result_wire[39] ;
wire \result_extra0_reg[39]~q ;
wire \result_wire[40] ;
wire \result_extra0_reg[40]~q ;
wire \result_wire[41] ;
wire \result_extra0_reg[41]~q ;
wire \result_wire[42] ;
wire \result_extra0_reg[42]~q ;
wire \result_wire[43] ;
wire \result_extra0_reg[43]~q ;
wire \result_wire[44] ;
wire \result_extra0_reg[44]~q ;
wire \result_wire[45] ;
wire \result_extra0_reg[45]~q ;
wire \result_wire[22] ;
wire \result_extra0_reg[22]~q ;
wire \result_wire[21] ;
wire \result_extra0_reg[21]~q ;
wire \result_wire[20] ;
wire \result_extra0_reg[20]~q ;
wire \result_wire[19] ;
wire \result_extra0_reg[19]~q ;
wire \result_wire[18] ;
wire \result_extra0_reg[18]~q ;
wire \result_wire[17] ;
wire \result_extra0_reg[17]~q ;
wire \result_wire[16] ;
wire \result_extra0_reg[16]~q ;
wire \result_wire[15] ;
wire \result_extra0_reg[15]~q ;
wire \result_wire[14] ;
wire \result_extra0_reg[14]~q ;
wire \result_wire[13] ;
wire \result_extra0_reg[13]~q ;
wire \result_wire[12] ;
wire \result_extra0_reg[12]~q ;
wire \result_wire[11] ;
wire \result_extra0_reg[11]~q ;
wire \result_wire[10] ;
wire \result_extra0_reg[10]~q ;
wire \result_wire[9] ;
wire \result_extra0_reg[9]~q ;
wire \result_wire[8] ;
wire \result_extra0_reg[8]~q ;
wire \result_wire[7] ;
wire \result_extra0_reg[7]~q ;
wire \result_wire[6] ;
wire \result_extra0_reg[6]~q ;
wire \result_wire[5] ;
wire \result_extra0_reg[5]~q ;
wire \result_wire[4] ;
wire \result_extra0_reg[4]~q ;
wire \result_wire[3] ;
wire \result_extra0_reg[3]~q ;
wire \result_wire[2] ;
wire \result_extra0_reg[2]~q ;
wire \result_wire[1] ;
wire \result_extra0_reg[1]~q ;
wire \result_wire[0] ;
wire \result_extra0_reg[0]~q ;

wire [63:0] \Mult0~mac_RESULTA_bus ;

assign \result_wire[0]  = \Mult0~mac_RESULTA_bus [0];
assign \result_wire[1]  = \Mult0~mac_RESULTA_bus [1];
assign \result_wire[2]  = \Mult0~mac_RESULTA_bus [2];
assign \result_wire[3]  = \Mult0~mac_RESULTA_bus [3];
assign \result_wire[4]  = \Mult0~mac_RESULTA_bus [4];
assign \result_wire[5]  = \Mult0~mac_RESULTA_bus [5];
assign \result_wire[6]  = \Mult0~mac_RESULTA_bus [6];
assign \result_wire[7]  = \Mult0~mac_RESULTA_bus [7];
assign \result_wire[8]  = \Mult0~mac_RESULTA_bus [8];
assign \result_wire[9]  = \Mult0~mac_RESULTA_bus [9];
assign \result_wire[10]  = \Mult0~mac_RESULTA_bus [10];
assign \result_wire[11]  = \Mult0~mac_RESULTA_bus [11];
assign \result_wire[12]  = \Mult0~mac_RESULTA_bus [12];
assign \result_wire[13]  = \Mult0~mac_RESULTA_bus [13];
assign \result_wire[14]  = \Mult0~mac_RESULTA_bus [14];
assign \result_wire[15]  = \Mult0~mac_RESULTA_bus [15];
assign \result_wire[16]  = \Mult0~mac_RESULTA_bus [16];
assign \result_wire[17]  = \Mult0~mac_RESULTA_bus [17];
assign \result_wire[18]  = \Mult0~mac_RESULTA_bus [18];
assign \result_wire[19]  = \Mult0~mac_RESULTA_bus [19];
assign \result_wire[20]  = \Mult0~mac_RESULTA_bus [20];
assign \result_wire[21]  = \Mult0~mac_RESULTA_bus [21];
assign \result_wire[22]  = \Mult0~mac_RESULTA_bus [22];
assign \result_wire[23]  = \Mult0~mac_RESULTA_bus [23];
assign \result_wire[24]  = \Mult0~mac_RESULTA_bus [24];
assign \result_wire[25]  = \Mult0~mac_RESULTA_bus [25];
assign \result_wire[26]  = \Mult0~mac_RESULTA_bus [26];
assign \result_wire[27]  = \Mult0~mac_RESULTA_bus [27];
assign \result_wire[28]  = \Mult0~mac_RESULTA_bus [28];
assign \result_wire[29]  = \Mult0~mac_RESULTA_bus [29];
assign \result_wire[30]  = \Mult0~mac_RESULTA_bus [30];
assign \result_wire[31]  = \Mult0~mac_RESULTA_bus [31];
assign \result_wire[32]  = \Mult0~mac_RESULTA_bus [32];
assign \result_wire[33]  = \Mult0~mac_RESULTA_bus [33];
assign \result_wire[34]  = \Mult0~mac_RESULTA_bus [34];
assign \result_wire[35]  = \Mult0~mac_RESULTA_bus [35];
assign \result_wire[36]  = \Mult0~mac_RESULTA_bus [36];
assign \result_wire[37]  = \Mult0~mac_RESULTA_bus [37];
assign \result_wire[38]  = \Mult0~mac_RESULTA_bus [38];
assign \result_wire[39]  = \Mult0~mac_RESULTA_bus [39];
assign \result_wire[40]  = \Mult0~mac_RESULTA_bus [40];
assign \result_wire[41]  = \Mult0~mac_RESULTA_bus [41];
assign \result_wire[42]  = \Mult0~mac_RESULTA_bus [42];
assign \result_wire[43]  = \Mult0~mac_RESULTA_bus [43];
assign \result_wire[44]  = \Mult0~mac_RESULTA_bus [44];
assign \result_wire[45]  = \Mult0~mac_RESULTA_bus [45];
assign \result_wire[46]  = \Mult0~mac_RESULTA_bus [46];
assign \result_wire[47]  = \Mult0~mac_RESULTA_bus [47];
assign \Mult0~8  = \Mult0~mac_RESULTA_bus [48];
assign \Mult0~9  = \Mult0~mac_RESULTA_bus [49];
assign \Mult0~10  = \Mult0~mac_RESULTA_bus [50];
assign \Mult0~11  = \Mult0~mac_RESULTA_bus [51];
assign \Mult0~12  = \Mult0~mac_RESULTA_bus [52];
assign \Mult0~13  = \Mult0~mac_RESULTA_bus [53];
assign \Mult0~14  = \Mult0~mac_RESULTA_bus [54];
assign \Mult0~15  = \Mult0~mac_RESULTA_bus [55];
assign \Mult0~16  = \Mult0~mac_RESULTA_bus [56];
assign \Mult0~17  = \Mult0~mac_RESULTA_bus [57];
assign \Mult0~18  = \Mult0~mac_RESULTA_bus [58];
assign \Mult0~19  = \Mult0~mac_RESULTA_bus [59];
assign \Mult0~20  = \Mult0~mac_RESULTA_bus [60];
assign \Mult0~21  = \Mult0~mac_RESULTA_bus [61];
assign \Mult0~22  = \Mult0~mac_RESULTA_bus [62];
assign \Mult0~23  = \Mult0~mac_RESULTA_bus [63];

dffeas \result_output_reg[46] (
	.clk(clock),
	.d(\result_extra0_reg[46]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_46),
	.prn(vcc));
defparam \result_output_reg[46] .is_wysiwyg = "true";
defparam \result_output_reg[46] .power_up = "low";

dffeas \result_output_reg[23] (
	.clk(clock),
	.d(\result_extra0_reg[23]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_23),
	.prn(vcc));
defparam \result_output_reg[23] .is_wysiwyg = "true";
defparam \result_output_reg[23] .power_up = "low";

dffeas \result_output_reg[34] (
	.clk(clock),
	.d(\result_extra0_reg[34]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_34),
	.prn(vcc));
defparam \result_output_reg[34] .is_wysiwyg = "true";
defparam \result_output_reg[34] .power_up = "low";

dffeas \result_output_reg[47] (
	.clk(clock),
	.d(\result_extra0_reg[47]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_47),
	.prn(vcc));
defparam \result_output_reg[47] .is_wysiwyg = "true";
defparam \result_output_reg[47] .power_up = "low";

dffeas \result_output_reg[24] (
	.clk(clock),
	.d(\result_extra0_reg[24]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_24),
	.prn(vcc));
defparam \result_output_reg[24] .is_wysiwyg = "true";
defparam \result_output_reg[24] .power_up = "low";

dffeas \result_output_reg[25] (
	.clk(clock),
	.d(\result_extra0_reg[25]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_25),
	.prn(vcc));
defparam \result_output_reg[25] .is_wysiwyg = "true";
defparam \result_output_reg[25] .power_up = "low";

dffeas \result_output_reg[26] (
	.clk(clock),
	.d(\result_extra0_reg[26]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_26),
	.prn(vcc));
defparam \result_output_reg[26] .is_wysiwyg = "true";
defparam \result_output_reg[26] .power_up = "low";

dffeas \result_output_reg[27] (
	.clk(clock),
	.d(\result_extra0_reg[27]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_27),
	.prn(vcc));
defparam \result_output_reg[27] .is_wysiwyg = "true";
defparam \result_output_reg[27] .power_up = "low";

dffeas \result_output_reg[28] (
	.clk(clock),
	.d(\result_extra0_reg[28]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_28),
	.prn(vcc));
defparam \result_output_reg[28] .is_wysiwyg = "true";
defparam \result_output_reg[28] .power_up = "low";

dffeas \result_output_reg[29] (
	.clk(clock),
	.d(\result_extra0_reg[29]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_29),
	.prn(vcc));
defparam \result_output_reg[29] .is_wysiwyg = "true";
defparam \result_output_reg[29] .power_up = "low";

dffeas \result_output_reg[30] (
	.clk(clock),
	.d(\result_extra0_reg[30]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_30),
	.prn(vcc));
defparam \result_output_reg[30] .is_wysiwyg = "true";
defparam \result_output_reg[30] .power_up = "low";

dffeas \result_output_reg[31] (
	.clk(clock),
	.d(\result_extra0_reg[31]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_31),
	.prn(vcc));
defparam \result_output_reg[31] .is_wysiwyg = "true";
defparam \result_output_reg[31] .power_up = "low";

dffeas \result_output_reg[32] (
	.clk(clock),
	.d(\result_extra0_reg[32]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_32),
	.prn(vcc));
defparam \result_output_reg[32] .is_wysiwyg = "true";
defparam \result_output_reg[32] .power_up = "low";

dffeas \result_output_reg[33] (
	.clk(clock),
	.d(\result_extra0_reg[33]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_33),
	.prn(vcc));
defparam \result_output_reg[33] .is_wysiwyg = "true";
defparam \result_output_reg[33] .power_up = "low";

dffeas \result_output_reg[35] (
	.clk(clock),
	.d(\result_extra0_reg[35]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_35),
	.prn(vcc));
defparam \result_output_reg[35] .is_wysiwyg = "true";
defparam \result_output_reg[35] .power_up = "low";

dffeas \result_output_reg[36] (
	.clk(clock),
	.d(\result_extra0_reg[36]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_36),
	.prn(vcc));
defparam \result_output_reg[36] .is_wysiwyg = "true";
defparam \result_output_reg[36] .power_up = "low";

dffeas \result_output_reg[37] (
	.clk(clock),
	.d(\result_extra0_reg[37]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_37),
	.prn(vcc));
defparam \result_output_reg[37] .is_wysiwyg = "true";
defparam \result_output_reg[37] .power_up = "low";

dffeas \result_output_reg[38] (
	.clk(clock),
	.d(\result_extra0_reg[38]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_38),
	.prn(vcc));
defparam \result_output_reg[38] .is_wysiwyg = "true";
defparam \result_output_reg[38] .power_up = "low";

dffeas \result_output_reg[39] (
	.clk(clock),
	.d(\result_extra0_reg[39]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_39),
	.prn(vcc));
defparam \result_output_reg[39] .is_wysiwyg = "true";
defparam \result_output_reg[39] .power_up = "low";

dffeas \result_output_reg[40] (
	.clk(clock),
	.d(\result_extra0_reg[40]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_40),
	.prn(vcc));
defparam \result_output_reg[40] .is_wysiwyg = "true";
defparam \result_output_reg[40] .power_up = "low";

dffeas \result_output_reg[41] (
	.clk(clock),
	.d(\result_extra0_reg[41]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_41),
	.prn(vcc));
defparam \result_output_reg[41] .is_wysiwyg = "true";
defparam \result_output_reg[41] .power_up = "low";

dffeas \result_output_reg[42] (
	.clk(clock),
	.d(\result_extra0_reg[42]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_42),
	.prn(vcc));
defparam \result_output_reg[42] .is_wysiwyg = "true";
defparam \result_output_reg[42] .power_up = "low";

dffeas \result_output_reg[43] (
	.clk(clock),
	.d(\result_extra0_reg[43]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_43),
	.prn(vcc));
defparam \result_output_reg[43] .is_wysiwyg = "true";
defparam \result_output_reg[43] .power_up = "low";

dffeas \result_output_reg[44] (
	.clk(clock),
	.d(\result_extra0_reg[44]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_44),
	.prn(vcc));
defparam \result_output_reg[44] .is_wysiwyg = "true";
defparam \result_output_reg[44] .power_up = "low";

dffeas \result_output_reg[45] (
	.clk(clock),
	.d(\result_extra0_reg[45]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_45),
	.prn(vcc));
defparam \result_output_reg[45] .is_wysiwyg = "true";
defparam \result_output_reg[45] .power_up = "low";

dffeas \result_output_reg[22] (
	.clk(clock),
	.d(\result_extra0_reg[22]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_22),
	.prn(vcc));
defparam \result_output_reg[22] .is_wysiwyg = "true";
defparam \result_output_reg[22] .power_up = "low";

dffeas \result_output_reg[21] (
	.clk(clock),
	.d(\result_extra0_reg[21]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_21),
	.prn(vcc));
defparam \result_output_reg[21] .is_wysiwyg = "true";
defparam \result_output_reg[21] .power_up = "low";

dffeas \result_output_reg[20] (
	.clk(clock),
	.d(\result_extra0_reg[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_20),
	.prn(vcc));
defparam \result_output_reg[20] .is_wysiwyg = "true";
defparam \result_output_reg[20] .power_up = "low";

dffeas \result_output_reg[19] (
	.clk(clock),
	.d(\result_extra0_reg[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_19),
	.prn(vcc));
defparam \result_output_reg[19] .is_wysiwyg = "true";
defparam \result_output_reg[19] .power_up = "low";

dffeas \result_output_reg[18] (
	.clk(clock),
	.d(\result_extra0_reg[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_18),
	.prn(vcc));
defparam \result_output_reg[18] .is_wysiwyg = "true";
defparam \result_output_reg[18] .power_up = "low";

dffeas \result_output_reg[17] (
	.clk(clock),
	.d(\result_extra0_reg[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_17),
	.prn(vcc));
defparam \result_output_reg[17] .is_wysiwyg = "true";
defparam \result_output_reg[17] .power_up = "low";

dffeas \result_output_reg[16] (
	.clk(clock),
	.d(\result_extra0_reg[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_16),
	.prn(vcc));
defparam \result_output_reg[16] .is_wysiwyg = "true";
defparam \result_output_reg[16] .power_up = "low";

dffeas \result_output_reg[15] (
	.clk(clock),
	.d(\result_extra0_reg[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_15),
	.prn(vcc));
defparam \result_output_reg[15] .is_wysiwyg = "true";
defparam \result_output_reg[15] .power_up = "low";

dffeas \result_output_reg[14] (
	.clk(clock),
	.d(\result_extra0_reg[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_14),
	.prn(vcc));
defparam \result_output_reg[14] .is_wysiwyg = "true";
defparam \result_output_reg[14] .power_up = "low";

dffeas \result_output_reg[13] (
	.clk(clock),
	.d(\result_extra0_reg[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_13),
	.prn(vcc));
defparam \result_output_reg[13] .is_wysiwyg = "true";
defparam \result_output_reg[13] .power_up = "low";

dffeas \result_output_reg[12] (
	.clk(clock),
	.d(\result_extra0_reg[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_12),
	.prn(vcc));
defparam \result_output_reg[12] .is_wysiwyg = "true";
defparam \result_output_reg[12] .power_up = "low";

dffeas \result_output_reg[11] (
	.clk(clock),
	.d(\result_extra0_reg[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_11),
	.prn(vcc));
defparam \result_output_reg[11] .is_wysiwyg = "true";
defparam \result_output_reg[11] .power_up = "low";

dffeas \result_output_reg[10] (
	.clk(clock),
	.d(\result_extra0_reg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_10),
	.prn(vcc));
defparam \result_output_reg[10] .is_wysiwyg = "true";
defparam \result_output_reg[10] .power_up = "low";

dffeas \result_output_reg[9] (
	.clk(clock),
	.d(\result_extra0_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_9),
	.prn(vcc));
defparam \result_output_reg[9] .is_wysiwyg = "true";
defparam \result_output_reg[9] .power_up = "low";

dffeas \result_output_reg[8] (
	.clk(clock),
	.d(\result_extra0_reg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_8),
	.prn(vcc));
defparam \result_output_reg[8] .is_wysiwyg = "true";
defparam \result_output_reg[8] .power_up = "low";

dffeas \result_output_reg[7] (
	.clk(clock),
	.d(\result_extra0_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_7),
	.prn(vcc));
defparam \result_output_reg[7] .is_wysiwyg = "true";
defparam \result_output_reg[7] .power_up = "low";

dffeas \result_output_reg[6] (
	.clk(clock),
	.d(\result_extra0_reg[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_6),
	.prn(vcc));
defparam \result_output_reg[6] .is_wysiwyg = "true";
defparam \result_output_reg[6] .power_up = "low";

dffeas \result_output_reg[5] (
	.clk(clock),
	.d(\result_extra0_reg[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_5),
	.prn(vcc));
defparam \result_output_reg[5] .is_wysiwyg = "true";
defparam \result_output_reg[5] .power_up = "low";

dffeas \result_output_reg[4] (
	.clk(clock),
	.d(\result_extra0_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_4),
	.prn(vcc));
defparam \result_output_reg[4] .is_wysiwyg = "true";
defparam \result_output_reg[4] .power_up = "low";

dffeas \result_output_reg[3] (
	.clk(clock),
	.d(\result_extra0_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_3),
	.prn(vcc));
defparam \result_output_reg[3] .is_wysiwyg = "true";
defparam \result_output_reg[3] .power_up = "low";

dffeas \result_output_reg[2] (
	.clk(clock),
	.d(\result_extra0_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_2),
	.prn(vcc));
defparam \result_output_reg[2] .is_wysiwyg = "true";
defparam \result_output_reg[2] .power_up = "low";

dffeas \result_output_reg[1] (
	.clk(clock),
	.d(\result_extra0_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_1),
	.prn(vcc));
defparam \result_output_reg[1] .is_wysiwyg = "true";
defparam \result_output_reg[1] .power_up = "low";

dffeas \result_output_reg[0] (
	.clk(clock),
	.d(\result_extra0_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_0),
	.prn(vcc));
defparam \result_output_reg[0] .is_wysiwyg = "true";
defparam \result_output_reg[0] .power_up = "low";

dffeas \dataa_input_reg[0] (
	.clk(clock),
	.d(dataa[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[0]~q ),
	.prn(vcc));
defparam \dataa_input_reg[0] .is_wysiwyg = "true";
defparam \dataa_input_reg[0] .power_up = "low";

dffeas \dataa_input_reg[1] (
	.clk(clock),
	.d(dataa[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[1]~q ),
	.prn(vcc));
defparam \dataa_input_reg[1] .is_wysiwyg = "true";
defparam \dataa_input_reg[1] .power_up = "low";

dffeas \dataa_input_reg[2] (
	.clk(clock),
	.d(dataa[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[2]~q ),
	.prn(vcc));
defparam \dataa_input_reg[2] .is_wysiwyg = "true";
defparam \dataa_input_reg[2] .power_up = "low";

dffeas \dataa_input_reg[3] (
	.clk(clock),
	.d(dataa[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[3]~q ),
	.prn(vcc));
defparam \dataa_input_reg[3] .is_wysiwyg = "true";
defparam \dataa_input_reg[3] .power_up = "low";

dffeas \dataa_input_reg[4] (
	.clk(clock),
	.d(dataa[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[4]~q ),
	.prn(vcc));
defparam \dataa_input_reg[4] .is_wysiwyg = "true";
defparam \dataa_input_reg[4] .power_up = "low";

dffeas \dataa_input_reg[5] (
	.clk(clock),
	.d(dataa[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[5]~q ),
	.prn(vcc));
defparam \dataa_input_reg[5] .is_wysiwyg = "true";
defparam \dataa_input_reg[5] .power_up = "low";

dffeas \dataa_input_reg[6] (
	.clk(clock),
	.d(dataa[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[6]~q ),
	.prn(vcc));
defparam \dataa_input_reg[6] .is_wysiwyg = "true";
defparam \dataa_input_reg[6] .power_up = "low";

dffeas \dataa_input_reg[7] (
	.clk(clock),
	.d(dataa[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[7]~q ),
	.prn(vcc));
defparam \dataa_input_reg[7] .is_wysiwyg = "true";
defparam \dataa_input_reg[7] .power_up = "low";

dffeas \dataa_input_reg[8] (
	.clk(clock),
	.d(dataa[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[8]~q ),
	.prn(vcc));
defparam \dataa_input_reg[8] .is_wysiwyg = "true";
defparam \dataa_input_reg[8] .power_up = "low";

dffeas \dataa_input_reg[9] (
	.clk(clock),
	.d(dataa[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[9]~q ),
	.prn(vcc));
defparam \dataa_input_reg[9] .is_wysiwyg = "true";
defparam \dataa_input_reg[9] .power_up = "low";

dffeas \dataa_input_reg[10] (
	.clk(clock),
	.d(dataa[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[10]~q ),
	.prn(vcc));
defparam \dataa_input_reg[10] .is_wysiwyg = "true";
defparam \dataa_input_reg[10] .power_up = "low";

dffeas \dataa_input_reg[11] (
	.clk(clock),
	.d(dataa[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[11]~q ),
	.prn(vcc));
defparam \dataa_input_reg[11] .is_wysiwyg = "true";
defparam \dataa_input_reg[11] .power_up = "low";

dffeas \dataa_input_reg[12] (
	.clk(clock),
	.d(dataa[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[12]~q ),
	.prn(vcc));
defparam \dataa_input_reg[12] .is_wysiwyg = "true";
defparam \dataa_input_reg[12] .power_up = "low";

dffeas \dataa_input_reg[13] (
	.clk(clock),
	.d(dataa[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[13]~q ),
	.prn(vcc));
defparam \dataa_input_reg[13] .is_wysiwyg = "true";
defparam \dataa_input_reg[13] .power_up = "low";

dffeas \dataa_input_reg[14] (
	.clk(clock),
	.d(dataa[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[14]~q ),
	.prn(vcc));
defparam \dataa_input_reg[14] .is_wysiwyg = "true";
defparam \dataa_input_reg[14] .power_up = "low";

dffeas \dataa_input_reg[15] (
	.clk(clock),
	.d(dataa[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[15]~q ),
	.prn(vcc));
defparam \dataa_input_reg[15] .is_wysiwyg = "true";
defparam \dataa_input_reg[15] .power_up = "low";

dffeas \dataa_input_reg[16] (
	.clk(clock),
	.d(dataa[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[16]~q ),
	.prn(vcc));
defparam \dataa_input_reg[16] .is_wysiwyg = "true";
defparam \dataa_input_reg[16] .power_up = "low";

dffeas \dataa_input_reg[17] (
	.clk(clock),
	.d(dataa[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[17]~q ),
	.prn(vcc));
defparam \dataa_input_reg[17] .is_wysiwyg = "true";
defparam \dataa_input_reg[17] .power_up = "low";

dffeas \dataa_input_reg[18] (
	.clk(clock),
	.d(dataa[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[18]~q ),
	.prn(vcc));
defparam \dataa_input_reg[18] .is_wysiwyg = "true";
defparam \dataa_input_reg[18] .power_up = "low";

dffeas \dataa_input_reg[19] (
	.clk(clock),
	.d(dataa[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[19]~q ),
	.prn(vcc));
defparam \dataa_input_reg[19] .is_wysiwyg = "true";
defparam \dataa_input_reg[19] .power_up = "low";

dffeas \dataa_input_reg[20] (
	.clk(clock),
	.d(dataa[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[20]~q ),
	.prn(vcc));
defparam \dataa_input_reg[20] .is_wysiwyg = "true";
defparam \dataa_input_reg[20] .power_up = "low";

dffeas \dataa_input_reg[21] (
	.clk(clock),
	.d(dataa[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[21]~q ),
	.prn(vcc));
defparam \dataa_input_reg[21] .is_wysiwyg = "true";
defparam \dataa_input_reg[21] .power_up = "low";

dffeas \dataa_input_reg[22] (
	.clk(clock),
	.d(dataa[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[22]~q ),
	.prn(vcc));
defparam \dataa_input_reg[22] .is_wysiwyg = "true";
defparam \dataa_input_reg[22] .power_up = "low";

dffeas \dataa_input_reg[23] (
	.clk(clock),
	.d(dataa[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[23]~q ),
	.prn(vcc));
defparam \dataa_input_reg[23] .is_wysiwyg = "true";
defparam \dataa_input_reg[23] .power_up = "low";

dffeas \datab_input_reg[0] (
	.clk(clock),
	.d(datab[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[0]~q ),
	.prn(vcc));
defparam \datab_input_reg[0] .is_wysiwyg = "true";
defparam \datab_input_reg[0] .power_up = "low";

dffeas \datab_input_reg[1] (
	.clk(clock),
	.d(datab[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[1]~q ),
	.prn(vcc));
defparam \datab_input_reg[1] .is_wysiwyg = "true";
defparam \datab_input_reg[1] .power_up = "low";

dffeas \datab_input_reg[2] (
	.clk(clock),
	.d(datab[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[2]~q ),
	.prn(vcc));
defparam \datab_input_reg[2] .is_wysiwyg = "true";
defparam \datab_input_reg[2] .power_up = "low";

dffeas \datab_input_reg[3] (
	.clk(clock),
	.d(datab[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[3]~q ),
	.prn(vcc));
defparam \datab_input_reg[3] .is_wysiwyg = "true";
defparam \datab_input_reg[3] .power_up = "low";

dffeas \datab_input_reg[4] (
	.clk(clock),
	.d(datab[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[4]~q ),
	.prn(vcc));
defparam \datab_input_reg[4] .is_wysiwyg = "true";
defparam \datab_input_reg[4] .power_up = "low";

dffeas \datab_input_reg[5] (
	.clk(clock),
	.d(datab[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[5]~q ),
	.prn(vcc));
defparam \datab_input_reg[5] .is_wysiwyg = "true";
defparam \datab_input_reg[5] .power_up = "low";

dffeas \datab_input_reg[6] (
	.clk(clock),
	.d(datab[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[6]~q ),
	.prn(vcc));
defparam \datab_input_reg[6] .is_wysiwyg = "true";
defparam \datab_input_reg[6] .power_up = "low";

dffeas \datab_input_reg[7] (
	.clk(clock),
	.d(datab[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[7]~q ),
	.prn(vcc));
defparam \datab_input_reg[7] .is_wysiwyg = "true";
defparam \datab_input_reg[7] .power_up = "low";

dffeas \datab_input_reg[8] (
	.clk(clock),
	.d(datab[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[8]~q ),
	.prn(vcc));
defparam \datab_input_reg[8] .is_wysiwyg = "true";
defparam \datab_input_reg[8] .power_up = "low";

dffeas \datab_input_reg[9] (
	.clk(clock),
	.d(datab[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[9]~q ),
	.prn(vcc));
defparam \datab_input_reg[9] .is_wysiwyg = "true";
defparam \datab_input_reg[9] .power_up = "low";

dffeas \datab_input_reg[10] (
	.clk(clock),
	.d(datab[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[10]~q ),
	.prn(vcc));
defparam \datab_input_reg[10] .is_wysiwyg = "true";
defparam \datab_input_reg[10] .power_up = "low";

dffeas \datab_input_reg[11] (
	.clk(clock),
	.d(datab[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[11]~q ),
	.prn(vcc));
defparam \datab_input_reg[11] .is_wysiwyg = "true";
defparam \datab_input_reg[11] .power_up = "low";

dffeas \datab_input_reg[12] (
	.clk(clock),
	.d(datab[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[12]~q ),
	.prn(vcc));
defparam \datab_input_reg[12] .is_wysiwyg = "true";
defparam \datab_input_reg[12] .power_up = "low";

dffeas \datab_input_reg[13] (
	.clk(clock),
	.d(datab[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[13]~q ),
	.prn(vcc));
defparam \datab_input_reg[13] .is_wysiwyg = "true";
defparam \datab_input_reg[13] .power_up = "low";

dffeas \datab_input_reg[14] (
	.clk(clock),
	.d(datab[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[14]~q ),
	.prn(vcc));
defparam \datab_input_reg[14] .is_wysiwyg = "true";
defparam \datab_input_reg[14] .power_up = "low";

dffeas \datab_input_reg[15] (
	.clk(clock),
	.d(datab[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[15]~q ),
	.prn(vcc));
defparam \datab_input_reg[15] .is_wysiwyg = "true";
defparam \datab_input_reg[15] .power_up = "low";

dffeas \datab_input_reg[16] (
	.clk(clock),
	.d(datab[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[16]~q ),
	.prn(vcc));
defparam \datab_input_reg[16] .is_wysiwyg = "true";
defparam \datab_input_reg[16] .power_up = "low";

dffeas \datab_input_reg[17] (
	.clk(clock),
	.d(datab[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[17]~q ),
	.prn(vcc));
defparam \datab_input_reg[17] .is_wysiwyg = "true";
defparam \datab_input_reg[17] .power_up = "low";

dffeas \datab_input_reg[18] (
	.clk(clock),
	.d(datab[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[18]~q ),
	.prn(vcc));
defparam \datab_input_reg[18] .is_wysiwyg = "true";
defparam \datab_input_reg[18] .power_up = "low";

dffeas \datab_input_reg[19] (
	.clk(clock),
	.d(datab[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[19]~q ),
	.prn(vcc));
defparam \datab_input_reg[19] .is_wysiwyg = "true";
defparam \datab_input_reg[19] .power_up = "low";

dffeas \datab_input_reg[20] (
	.clk(clock),
	.d(datab[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[20]~q ),
	.prn(vcc));
defparam \datab_input_reg[20] .is_wysiwyg = "true";
defparam \datab_input_reg[20] .power_up = "low";

dffeas \datab_input_reg[21] (
	.clk(clock),
	.d(datab[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[21]~q ),
	.prn(vcc));
defparam \datab_input_reg[21] .is_wysiwyg = "true";
defparam \datab_input_reg[21] .power_up = "low";

dffeas \datab_input_reg[22] (
	.clk(clock),
	.d(datab[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[22]~q ),
	.prn(vcc));
defparam \datab_input_reg[22] .is_wysiwyg = "true";
defparam \datab_input_reg[22] .power_up = "low";

dffeas \datab_input_reg[23] (
	.clk(clock),
	.d(datab[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[23]~q ),
	.prn(vcc));
defparam \datab_input_reg[23] .is_wysiwyg = "true";
defparam \datab_input_reg[23] .power_up = "low";

cyclonev_mac \Mult0~mac (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,\dataa_input_reg[23]~q ,\dataa_input_reg[22]~q ,\dataa_input_reg[21]~q ,\dataa_input_reg[20]~q ,\dataa_input_reg[19]~q ,\dataa_input_reg[18]~q ,\dataa_input_reg[17]~q ,\dataa_input_reg[16]~q ,\dataa_input_reg[15]~q ,\dataa_input_reg[14]~q ,
\dataa_input_reg[13]~q ,\dataa_input_reg[12]~q ,\dataa_input_reg[11]~q ,\dataa_input_reg[10]~q ,\dataa_input_reg[9]~q ,\dataa_input_reg[8]~q ,\dataa_input_reg[7]~q ,\dataa_input_reg[6]~q ,\dataa_input_reg[5]~q ,\dataa_input_reg[4]~q ,\dataa_input_reg[3]~q ,
\dataa_input_reg[2]~q ,\dataa_input_reg[1]~q ,\dataa_input_reg[0]~q }),
	.ay({gnd,gnd,gnd,\datab_input_reg[23]~q ,\datab_input_reg[22]~q ,\datab_input_reg[21]~q ,\datab_input_reg[20]~q ,\datab_input_reg[19]~q ,\datab_input_reg[18]~q ,\datab_input_reg[17]~q ,\datab_input_reg[16]~q ,\datab_input_reg[15]~q ,\datab_input_reg[14]~q ,
\datab_input_reg[13]~q ,\datab_input_reg[12]~q ,\datab_input_reg[11]~q ,\datab_input_reg[10]~q ,\datab_input_reg[9]~q ,\datab_input_reg[8]~q ,\datab_input_reg[7]~q ,\datab_input_reg[6]~q ,\datab_input_reg[5]~q ,\datab_input_reg[4]~q ,\datab_input_reg[3]~q ,
\datab_input_reg[2]~q ,\datab_input_reg[1]~q ,\datab_input_reg[0]~q }),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Mult0~mac_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Mult0~mac .accumulate_clock = "none";
defparam \Mult0~mac .ax_clock = "none";
defparam \Mult0~mac .ax_width = 24;
defparam \Mult0~mac .ay_scan_in_clock = "none";
defparam \Mult0~mac .ay_scan_in_width = 24;
defparam \Mult0~mac .ay_use_scan_in = "false";
defparam \Mult0~mac .az_clock = "none";
defparam \Mult0~mac .bx_clock = "none";
defparam \Mult0~mac .by_clock = "none";
defparam \Mult0~mac .by_use_scan_in = "false";
defparam \Mult0~mac .bz_clock = "none";
defparam \Mult0~mac .coef_a_0 = 0;
defparam \Mult0~mac .coef_a_1 = 0;
defparam \Mult0~mac .coef_a_2 = 0;
defparam \Mult0~mac .coef_a_3 = 0;
defparam \Mult0~mac .coef_a_4 = 0;
defparam \Mult0~mac .coef_a_5 = 0;
defparam \Mult0~mac .coef_a_6 = 0;
defparam \Mult0~mac .coef_a_7 = 0;
defparam \Mult0~mac .coef_b_0 = 0;
defparam \Mult0~mac .coef_b_1 = 0;
defparam \Mult0~mac .coef_b_2 = 0;
defparam \Mult0~mac .coef_b_3 = 0;
defparam \Mult0~mac .coef_b_4 = 0;
defparam \Mult0~mac .coef_b_5 = 0;
defparam \Mult0~mac .coef_b_6 = 0;
defparam \Mult0~mac .coef_b_7 = 0;
defparam \Mult0~mac .coef_sel_a_clock = "none";
defparam \Mult0~mac .coef_sel_b_clock = "none";
defparam \Mult0~mac .delay_scan_out_ay = "false";
defparam \Mult0~mac .delay_scan_out_by = "false";
defparam \Mult0~mac .enable_double_accum = "false";
defparam \Mult0~mac .load_const_clock = "none";
defparam \Mult0~mac .load_const_value = 0;
defparam \Mult0~mac .mode_sub_location = 0;
defparam \Mult0~mac .negate_clock = "none";
defparam \Mult0~mac .operand_source_max = "input";
defparam \Mult0~mac .operand_source_may = "input";
defparam \Mult0~mac .operand_source_mbx = "input";
defparam \Mult0~mac .operand_source_mby = "input";
defparam \Mult0~mac .operation_mode = "m27x27";
defparam \Mult0~mac .output_clock = "none";
defparam \Mult0~mac .preadder_subtract_a = "false";
defparam \Mult0~mac .preadder_subtract_b = "false";
defparam \Mult0~mac .result_a_width = 64;
defparam \Mult0~mac .signed_max = "true";
defparam \Mult0~mac .signed_may = "true";
defparam \Mult0~mac .signed_mbx = "false";
defparam \Mult0~mac .signed_mby = "false";
defparam \Mult0~mac .sub_clock = "none";
defparam \Mult0~mac .use_chainadder = "false";

dffeas \result_extra0_reg[46] (
	.clk(clock),
	.d(\result_wire[46] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[46]~q ),
	.prn(vcc));
defparam \result_extra0_reg[46] .is_wysiwyg = "true";
defparam \result_extra0_reg[46] .power_up = "low";

dffeas \result_extra0_reg[23] (
	.clk(clock),
	.d(\result_wire[23] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[23]~q ),
	.prn(vcc));
defparam \result_extra0_reg[23] .is_wysiwyg = "true";
defparam \result_extra0_reg[23] .power_up = "low";

dffeas \result_extra0_reg[34] (
	.clk(clock),
	.d(\result_wire[34] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[34]~q ),
	.prn(vcc));
defparam \result_extra0_reg[34] .is_wysiwyg = "true";
defparam \result_extra0_reg[34] .power_up = "low";

dffeas \result_extra0_reg[47] (
	.clk(clock),
	.d(\result_wire[47] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[47]~q ),
	.prn(vcc));
defparam \result_extra0_reg[47] .is_wysiwyg = "true";
defparam \result_extra0_reg[47] .power_up = "low";

dffeas \result_extra0_reg[24] (
	.clk(clock),
	.d(\result_wire[24] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[24]~q ),
	.prn(vcc));
defparam \result_extra0_reg[24] .is_wysiwyg = "true";
defparam \result_extra0_reg[24] .power_up = "low";

dffeas \result_extra0_reg[25] (
	.clk(clock),
	.d(\result_wire[25] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[25]~q ),
	.prn(vcc));
defparam \result_extra0_reg[25] .is_wysiwyg = "true";
defparam \result_extra0_reg[25] .power_up = "low";

dffeas \result_extra0_reg[26] (
	.clk(clock),
	.d(\result_wire[26] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[26]~q ),
	.prn(vcc));
defparam \result_extra0_reg[26] .is_wysiwyg = "true";
defparam \result_extra0_reg[26] .power_up = "low";

dffeas \result_extra0_reg[27] (
	.clk(clock),
	.d(\result_wire[27] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[27]~q ),
	.prn(vcc));
defparam \result_extra0_reg[27] .is_wysiwyg = "true";
defparam \result_extra0_reg[27] .power_up = "low";

dffeas \result_extra0_reg[28] (
	.clk(clock),
	.d(\result_wire[28] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[28]~q ),
	.prn(vcc));
defparam \result_extra0_reg[28] .is_wysiwyg = "true";
defparam \result_extra0_reg[28] .power_up = "low";

dffeas \result_extra0_reg[29] (
	.clk(clock),
	.d(\result_wire[29] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[29]~q ),
	.prn(vcc));
defparam \result_extra0_reg[29] .is_wysiwyg = "true";
defparam \result_extra0_reg[29] .power_up = "low";

dffeas \result_extra0_reg[30] (
	.clk(clock),
	.d(\result_wire[30] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[30]~q ),
	.prn(vcc));
defparam \result_extra0_reg[30] .is_wysiwyg = "true";
defparam \result_extra0_reg[30] .power_up = "low";

dffeas \result_extra0_reg[31] (
	.clk(clock),
	.d(\result_wire[31] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[31]~q ),
	.prn(vcc));
defparam \result_extra0_reg[31] .is_wysiwyg = "true";
defparam \result_extra0_reg[31] .power_up = "low";

dffeas \result_extra0_reg[32] (
	.clk(clock),
	.d(\result_wire[32] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[32]~q ),
	.prn(vcc));
defparam \result_extra0_reg[32] .is_wysiwyg = "true";
defparam \result_extra0_reg[32] .power_up = "low";

dffeas \result_extra0_reg[33] (
	.clk(clock),
	.d(\result_wire[33] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[33]~q ),
	.prn(vcc));
defparam \result_extra0_reg[33] .is_wysiwyg = "true";
defparam \result_extra0_reg[33] .power_up = "low";

dffeas \result_extra0_reg[35] (
	.clk(clock),
	.d(\result_wire[35] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[35]~q ),
	.prn(vcc));
defparam \result_extra0_reg[35] .is_wysiwyg = "true";
defparam \result_extra0_reg[35] .power_up = "low";

dffeas \result_extra0_reg[36] (
	.clk(clock),
	.d(\result_wire[36] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[36]~q ),
	.prn(vcc));
defparam \result_extra0_reg[36] .is_wysiwyg = "true";
defparam \result_extra0_reg[36] .power_up = "low";

dffeas \result_extra0_reg[37] (
	.clk(clock),
	.d(\result_wire[37] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[37]~q ),
	.prn(vcc));
defparam \result_extra0_reg[37] .is_wysiwyg = "true";
defparam \result_extra0_reg[37] .power_up = "low";

dffeas \result_extra0_reg[38] (
	.clk(clock),
	.d(\result_wire[38] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[38]~q ),
	.prn(vcc));
defparam \result_extra0_reg[38] .is_wysiwyg = "true";
defparam \result_extra0_reg[38] .power_up = "low";

dffeas \result_extra0_reg[39] (
	.clk(clock),
	.d(\result_wire[39] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[39]~q ),
	.prn(vcc));
defparam \result_extra0_reg[39] .is_wysiwyg = "true";
defparam \result_extra0_reg[39] .power_up = "low";

dffeas \result_extra0_reg[40] (
	.clk(clock),
	.d(\result_wire[40] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[40]~q ),
	.prn(vcc));
defparam \result_extra0_reg[40] .is_wysiwyg = "true";
defparam \result_extra0_reg[40] .power_up = "low";

dffeas \result_extra0_reg[41] (
	.clk(clock),
	.d(\result_wire[41] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[41]~q ),
	.prn(vcc));
defparam \result_extra0_reg[41] .is_wysiwyg = "true";
defparam \result_extra0_reg[41] .power_up = "low";

dffeas \result_extra0_reg[42] (
	.clk(clock),
	.d(\result_wire[42] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[42]~q ),
	.prn(vcc));
defparam \result_extra0_reg[42] .is_wysiwyg = "true";
defparam \result_extra0_reg[42] .power_up = "low";

dffeas \result_extra0_reg[43] (
	.clk(clock),
	.d(\result_wire[43] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[43]~q ),
	.prn(vcc));
defparam \result_extra0_reg[43] .is_wysiwyg = "true";
defparam \result_extra0_reg[43] .power_up = "low";

dffeas \result_extra0_reg[44] (
	.clk(clock),
	.d(\result_wire[44] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[44]~q ),
	.prn(vcc));
defparam \result_extra0_reg[44] .is_wysiwyg = "true";
defparam \result_extra0_reg[44] .power_up = "low";

dffeas \result_extra0_reg[45] (
	.clk(clock),
	.d(\result_wire[45] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[45]~q ),
	.prn(vcc));
defparam \result_extra0_reg[45] .is_wysiwyg = "true";
defparam \result_extra0_reg[45] .power_up = "low";

dffeas \result_extra0_reg[22] (
	.clk(clock),
	.d(\result_wire[22] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[22]~q ),
	.prn(vcc));
defparam \result_extra0_reg[22] .is_wysiwyg = "true";
defparam \result_extra0_reg[22] .power_up = "low";

dffeas \result_extra0_reg[21] (
	.clk(clock),
	.d(\result_wire[21] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[21]~q ),
	.prn(vcc));
defparam \result_extra0_reg[21] .is_wysiwyg = "true";
defparam \result_extra0_reg[21] .power_up = "low";

dffeas \result_extra0_reg[20] (
	.clk(clock),
	.d(\result_wire[20] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[20]~q ),
	.prn(vcc));
defparam \result_extra0_reg[20] .is_wysiwyg = "true";
defparam \result_extra0_reg[20] .power_up = "low";

dffeas \result_extra0_reg[19] (
	.clk(clock),
	.d(\result_wire[19] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[19]~q ),
	.prn(vcc));
defparam \result_extra0_reg[19] .is_wysiwyg = "true";
defparam \result_extra0_reg[19] .power_up = "low";

dffeas \result_extra0_reg[18] (
	.clk(clock),
	.d(\result_wire[18] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[18]~q ),
	.prn(vcc));
defparam \result_extra0_reg[18] .is_wysiwyg = "true";
defparam \result_extra0_reg[18] .power_up = "low";

dffeas \result_extra0_reg[17] (
	.clk(clock),
	.d(\result_wire[17] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[17]~q ),
	.prn(vcc));
defparam \result_extra0_reg[17] .is_wysiwyg = "true";
defparam \result_extra0_reg[17] .power_up = "low";

dffeas \result_extra0_reg[16] (
	.clk(clock),
	.d(\result_wire[16] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[16]~q ),
	.prn(vcc));
defparam \result_extra0_reg[16] .is_wysiwyg = "true";
defparam \result_extra0_reg[16] .power_up = "low";

dffeas \result_extra0_reg[15] (
	.clk(clock),
	.d(\result_wire[15] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[15]~q ),
	.prn(vcc));
defparam \result_extra0_reg[15] .is_wysiwyg = "true";
defparam \result_extra0_reg[15] .power_up = "low";

dffeas \result_extra0_reg[14] (
	.clk(clock),
	.d(\result_wire[14] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[14]~q ),
	.prn(vcc));
defparam \result_extra0_reg[14] .is_wysiwyg = "true";
defparam \result_extra0_reg[14] .power_up = "low";

dffeas \result_extra0_reg[13] (
	.clk(clock),
	.d(\result_wire[13] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[13]~q ),
	.prn(vcc));
defparam \result_extra0_reg[13] .is_wysiwyg = "true";
defparam \result_extra0_reg[13] .power_up = "low";

dffeas \result_extra0_reg[12] (
	.clk(clock),
	.d(\result_wire[12] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[12]~q ),
	.prn(vcc));
defparam \result_extra0_reg[12] .is_wysiwyg = "true";
defparam \result_extra0_reg[12] .power_up = "low";

dffeas \result_extra0_reg[11] (
	.clk(clock),
	.d(\result_wire[11] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[11]~q ),
	.prn(vcc));
defparam \result_extra0_reg[11] .is_wysiwyg = "true";
defparam \result_extra0_reg[11] .power_up = "low";

dffeas \result_extra0_reg[10] (
	.clk(clock),
	.d(\result_wire[10] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[10]~q ),
	.prn(vcc));
defparam \result_extra0_reg[10] .is_wysiwyg = "true";
defparam \result_extra0_reg[10] .power_up = "low";

dffeas \result_extra0_reg[9] (
	.clk(clock),
	.d(\result_wire[9] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[9]~q ),
	.prn(vcc));
defparam \result_extra0_reg[9] .is_wysiwyg = "true";
defparam \result_extra0_reg[9] .power_up = "low";

dffeas \result_extra0_reg[8] (
	.clk(clock),
	.d(\result_wire[8] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[8]~q ),
	.prn(vcc));
defparam \result_extra0_reg[8] .is_wysiwyg = "true";
defparam \result_extra0_reg[8] .power_up = "low";

dffeas \result_extra0_reg[7] (
	.clk(clock),
	.d(\result_wire[7] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[7]~q ),
	.prn(vcc));
defparam \result_extra0_reg[7] .is_wysiwyg = "true";
defparam \result_extra0_reg[7] .power_up = "low";

dffeas \result_extra0_reg[6] (
	.clk(clock),
	.d(\result_wire[6] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[6]~q ),
	.prn(vcc));
defparam \result_extra0_reg[6] .is_wysiwyg = "true";
defparam \result_extra0_reg[6] .power_up = "low";

dffeas \result_extra0_reg[5] (
	.clk(clock),
	.d(\result_wire[5] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[5]~q ),
	.prn(vcc));
defparam \result_extra0_reg[5] .is_wysiwyg = "true";
defparam \result_extra0_reg[5] .power_up = "low";

dffeas \result_extra0_reg[4] (
	.clk(clock),
	.d(\result_wire[4] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[4]~q ),
	.prn(vcc));
defparam \result_extra0_reg[4] .is_wysiwyg = "true";
defparam \result_extra0_reg[4] .power_up = "low";

dffeas \result_extra0_reg[3] (
	.clk(clock),
	.d(\result_wire[3] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[3]~q ),
	.prn(vcc));
defparam \result_extra0_reg[3] .is_wysiwyg = "true";
defparam \result_extra0_reg[3] .power_up = "low";

dffeas \result_extra0_reg[2] (
	.clk(clock),
	.d(\result_wire[2] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[2]~q ),
	.prn(vcc));
defparam \result_extra0_reg[2] .is_wysiwyg = "true";
defparam \result_extra0_reg[2] .power_up = "low";

dffeas \result_extra0_reg[1] (
	.clk(clock),
	.d(\result_wire[1] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[1]~q ),
	.prn(vcc));
defparam \result_extra0_reg[1] .is_wysiwyg = "true";
defparam \result_extra0_reg[1] .power_up = "low";

dffeas \result_extra0_reg[0] (
	.clk(clock),
	.d(\result_wire[0] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[0]~q ),
	.prn(vcc));
defparam \result_extra0_reg[0] .is_wysiwyg = "true";
defparam \result_extra0_reg[0] .power_up = "low";

endmodule

module sine_lmsd_1 (
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_21,
	q_b_22,
	q_b_23,
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_8,
	q_a_9,
	q_a_10,
	q_a_11,
	q_a_12,
	q_a_13,
	q_a_14,
	q_a_15,
	q_a_16,
	q_a_17,
	q_a_18,
	q_a_19,
	q_a_20,
	q_a_21,
	q_a_22,
	q_a_23,
	result_output_reg_46,
	result_output_reg_23,
	result_output_reg_34,
	result_output_reg_47,
	result_output_reg_24,
	result_output_reg_25,
	result_output_reg_26,
	result_output_reg_27,
	result_output_reg_28,
	result_output_reg_29,
	result_output_reg_30,
	result_output_reg_31,
	result_output_reg_32,
	result_output_reg_33,
	result_output_reg_35,
	result_output_reg_36,
	result_output_reg_37,
	result_output_reg_38,
	result_output_reg_39,
	result_output_reg_40,
	result_output_reg_41,
	result_output_reg_42,
	result_output_reg_43,
	result_output_reg_44,
	result_output_reg_45,
	result_output_reg_22,
	result_output_reg_21,
	result_output_reg_20,
	result_output_reg_19,
	result_output_reg_18,
	result_output_reg_17,
	result_output_reg_16,
	result_output_reg_15,
	result_output_reg_14,
	result_output_reg_13,
	result_output_reg_12,
	result_output_reg_11,
	result_output_reg_10,
	result_output_reg_9,
	result_output_reg_8,
	result_output_reg_7,
	result_output_reg_6,
	result_output_reg_5,
	result_output_reg_4,
	result_output_reg_3,
	result_output_reg_2,
	result_output_reg_1,
	result_output_reg_0,
	clk,
	clken)/* synthesis synthesis_greybox=1 */;
input 	q_b_0;
input 	q_b_1;
input 	q_b_2;
input 	q_b_3;
input 	q_b_4;
input 	q_b_5;
input 	q_b_6;
input 	q_b_7;
input 	q_b_8;
input 	q_b_9;
input 	q_b_10;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_20;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_a_0;
input 	q_a_1;
input 	q_a_2;
input 	q_a_3;
input 	q_a_4;
input 	q_a_5;
input 	q_a_6;
input 	q_a_7;
input 	q_a_8;
input 	q_a_9;
input 	q_a_10;
input 	q_a_11;
input 	q_a_12;
input 	q_a_13;
input 	q_a_14;
input 	q_a_15;
input 	q_a_16;
input 	q_a_17;
input 	q_a_18;
input 	q_a_19;
input 	q_a_20;
input 	q_a_21;
input 	q_a_22;
input 	q_a_23;
output 	result_output_reg_46;
output 	result_output_reg_23;
output 	result_output_reg_34;
output 	result_output_reg_47;
output 	result_output_reg_24;
output 	result_output_reg_25;
output 	result_output_reg_26;
output 	result_output_reg_27;
output 	result_output_reg_28;
output 	result_output_reg_29;
output 	result_output_reg_30;
output 	result_output_reg_31;
output 	result_output_reg_32;
output 	result_output_reg_33;
output 	result_output_reg_35;
output 	result_output_reg_36;
output 	result_output_reg_37;
output 	result_output_reg_38;
output 	result_output_reg_39;
output 	result_output_reg_40;
output 	result_output_reg_41;
output 	result_output_reg_42;
output 	result_output_reg_43;
output 	result_output_reg_44;
output 	result_output_reg_45;
output 	result_output_reg_22;
output 	result_output_reg_21;
output 	result_output_reg_20;
output 	result_output_reg_19;
output 	result_output_reg_18;
output 	result_output_reg_17;
output 	result_output_reg_16;
output 	result_output_reg_15;
output 	result_output_reg_14;
output 	result_output_reg_13;
output 	result_output_reg_12;
output 	result_output_reg_11;
output 	result_output_reg_10;
output 	result_output_reg_9;
output 	result_output_reg_8;
output 	result_output_reg_7;
output 	result_output_reg_6;
output 	result_output_reg_5;
output 	result_output_reg_4;
output 	result_output_reg_3;
output 	result_output_reg_2;
output 	result_output_reg_1;
output 	result_output_reg_0;
input 	clk;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_lpm_mult_2 lpm_mult_component(
	.datab({q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.dataa({q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.result_output_reg_46(result_output_reg_46),
	.result_output_reg_23(result_output_reg_23),
	.result_output_reg_34(result_output_reg_34),
	.result_output_reg_47(result_output_reg_47),
	.result_output_reg_24(result_output_reg_24),
	.result_output_reg_25(result_output_reg_25),
	.result_output_reg_26(result_output_reg_26),
	.result_output_reg_27(result_output_reg_27),
	.result_output_reg_28(result_output_reg_28),
	.result_output_reg_29(result_output_reg_29),
	.result_output_reg_30(result_output_reg_30),
	.result_output_reg_31(result_output_reg_31),
	.result_output_reg_32(result_output_reg_32),
	.result_output_reg_33(result_output_reg_33),
	.result_output_reg_35(result_output_reg_35),
	.result_output_reg_36(result_output_reg_36),
	.result_output_reg_37(result_output_reg_37),
	.result_output_reg_38(result_output_reg_38),
	.result_output_reg_39(result_output_reg_39),
	.result_output_reg_40(result_output_reg_40),
	.result_output_reg_41(result_output_reg_41),
	.result_output_reg_42(result_output_reg_42),
	.result_output_reg_43(result_output_reg_43),
	.result_output_reg_44(result_output_reg_44),
	.result_output_reg_45(result_output_reg_45),
	.result_output_reg_22(result_output_reg_22),
	.result_output_reg_21(result_output_reg_21),
	.result_output_reg_20(result_output_reg_20),
	.result_output_reg_19(result_output_reg_19),
	.result_output_reg_18(result_output_reg_18),
	.result_output_reg_17(result_output_reg_17),
	.result_output_reg_16(result_output_reg_16),
	.result_output_reg_15(result_output_reg_15),
	.result_output_reg_14(result_output_reg_14),
	.result_output_reg_13(result_output_reg_13),
	.result_output_reg_12(result_output_reg_12),
	.result_output_reg_11(result_output_reg_11),
	.result_output_reg_10(result_output_reg_10),
	.result_output_reg_9(result_output_reg_9),
	.result_output_reg_8(result_output_reg_8),
	.result_output_reg_7(result_output_reg_7),
	.result_output_reg_6(result_output_reg_6),
	.result_output_reg_5(result_output_reg_5),
	.result_output_reg_4(result_output_reg_4),
	.result_output_reg_3(result_output_reg_3),
	.result_output_reg_2(result_output_reg_2),
	.result_output_reg_1(result_output_reg_1),
	.result_output_reg_0(result_output_reg_0),
	.clock(clk),
	.clken(clken));

endmodule

module sine_lpm_mult_2 (
	datab,
	dataa,
	result_output_reg_46,
	result_output_reg_23,
	result_output_reg_34,
	result_output_reg_47,
	result_output_reg_24,
	result_output_reg_25,
	result_output_reg_26,
	result_output_reg_27,
	result_output_reg_28,
	result_output_reg_29,
	result_output_reg_30,
	result_output_reg_31,
	result_output_reg_32,
	result_output_reg_33,
	result_output_reg_35,
	result_output_reg_36,
	result_output_reg_37,
	result_output_reg_38,
	result_output_reg_39,
	result_output_reg_40,
	result_output_reg_41,
	result_output_reg_42,
	result_output_reg_43,
	result_output_reg_44,
	result_output_reg_45,
	result_output_reg_22,
	result_output_reg_21,
	result_output_reg_20,
	result_output_reg_19,
	result_output_reg_18,
	result_output_reg_17,
	result_output_reg_16,
	result_output_reg_15,
	result_output_reg_14,
	result_output_reg_13,
	result_output_reg_12,
	result_output_reg_11,
	result_output_reg_10,
	result_output_reg_9,
	result_output_reg_8,
	result_output_reg_7,
	result_output_reg_6,
	result_output_reg_5,
	result_output_reg_4,
	result_output_reg_3,
	result_output_reg_2,
	result_output_reg_1,
	result_output_reg_0,
	clock,
	clken)/* synthesis synthesis_greybox=1 */;
input 	[23:0] datab;
input 	[23:0] dataa;
output 	result_output_reg_46;
output 	result_output_reg_23;
output 	result_output_reg_34;
output 	result_output_reg_47;
output 	result_output_reg_24;
output 	result_output_reg_25;
output 	result_output_reg_26;
output 	result_output_reg_27;
output 	result_output_reg_28;
output 	result_output_reg_29;
output 	result_output_reg_30;
output 	result_output_reg_31;
output 	result_output_reg_32;
output 	result_output_reg_33;
output 	result_output_reg_35;
output 	result_output_reg_36;
output 	result_output_reg_37;
output 	result_output_reg_38;
output 	result_output_reg_39;
output 	result_output_reg_40;
output 	result_output_reg_41;
output 	result_output_reg_42;
output 	result_output_reg_43;
output 	result_output_reg_44;
output 	result_output_reg_45;
output 	result_output_reg_22;
output 	result_output_reg_21;
output 	result_output_reg_20;
output 	result_output_reg_19;
output 	result_output_reg_18;
output 	result_output_reg_17;
output 	result_output_reg_16;
output 	result_output_reg_15;
output 	result_output_reg_14;
output 	result_output_reg_13;
output 	result_output_reg_12;
output 	result_output_reg_11;
output 	result_output_reg_10;
output 	result_output_reg_9;
output 	result_output_reg_8;
output 	result_output_reg_7;
output 	result_output_reg_6;
output 	result_output_reg_5;
output 	result_output_reg_4;
output 	result_output_reg_3;
output 	result_output_reg_2;
output 	result_output_reg_1;
output 	result_output_reg_0;
input 	clock;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_mult_5cu_1 auto_generated(
	.datab({datab[23],datab[22],datab[21],datab[20],datab[19],datab[18],datab[17],datab[16],datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataa({dataa[23],dataa[22],dataa[21],dataa[20],dataa[19],dataa[18],dataa[17],dataa[16],dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.result_output_reg_46(result_output_reg_46),
	.result_output_reg_23(result_output_reg_23),
	.result_output_reg_34(result_output_reg_34),
	.result_output_reg_47(result_output_reg_47),
	.result_output_reg_24(result_output_reg_24),
	.result_output_reg_25(result_output_reg_25),
	.result_output_reg_26(result_output_reg_26),
	.result_output_reg_27(result_output_reg_27),
	.result_output_reg_28(result_output_reg_28),
	.result_output_reg_29(result_output_reg_29),
	.result_output_reg_30(result_output_reg_30),
	.result_output_reg_31(result_output_reg_31),
	.result_output_reg_32(result_output_reg_32),
	.result_output_reg_33(result_output_reg_33),
	.result_output_reg_35(result_output_reg_35),
	.result_output_reg_36(result_output_reg_36),
	.result_output_reg_37(result_output_reg_37),
	.result_output_reg_38(result_output_reg_38),
	.result_output_reg_39(result_output_reg_39),
	.result_output_reg_40(result_output_reg_40),
	.result_output_reg_41(result_output_reg_41),
	.result_output_reg_42(result_output_reg_42),
	.result_output_reg_43(result_output_reg_43),
	.result_output_reg_44(result_output_reg_44),
	.result_output_reg_45(result_output_reg_45),
	.result_output_reg_22(result_output_reg_22),
	.result_output_reg_21(result_output_reg_21),
	.result_output_reg_20(result_output_reg_20),
	.result_output_reg_19(result_output_reg_19),
	.result_output_reg_18(result_output_reg_18),
	.result_output_reg_17(result_output_reg_17),
	.result_output_reg_16(result_output_reg_16),
	.result_output_reg_15(result_output_reg_15),
	.result_output_reg_14(result_output_reg_14),
	.result_output_reg_13(result_output_reg_13),
	.result_output_reg_12(result_output_reg_12),
	.result_output_reg_11(result_output_reg_11),
	.result_output_reg_10(result_output_reg_10),
	.result_output_reg_9(result_output_reg_9),
	.result_output_reg_8(result_output_reg_8),
	.result_output_reg_7(result_output_reg_7),
	.result_output_reg_6(result_output_reg_6),
	.result_output_reg_5(result_output_reg_5),
	.result_output_reg_4(result_output_reg_4),
	.result_output_reg_3(result_output_reg_3),
	.result_output_reg_2(result_output_reg_2),
	.result_output_reg_1(result_output_reg_1),
	.result_output_reg_0(result_output_reg_0),
	.clock(clock),
	.clken(clken));

endmodule

module sine_mult_5cu_1 (
	datab,
	dataa,
	result_output_reg_46,
	result_output_reg_23,
	result_output_reg_34,
	result_output_reg_47,
	result_output_reg_24,
	result_output_reg_25,
	result_output_reg_26,
	result_output_reg_27,
	result_output_reg_28,
	result_output_reg_29,
	result_output_reg_30,
	result_output_reg_31,
	result_output_reg_32,
	result_output_reg_33,
	result_output_reg_35,
	result_output_reg_36,
	result_output_reg_37,
	result_output_reg_38,
	result_output_reg_39,
	result_output_reg_40,
	result_output_reg_41,
	result_output_reg_42,
	result_output_reg_43,
	result_output_reg_44,
	result_output_reg_45,
	result_output_reg_22,
	result_output_reg_21,
	result_output_reg_20,
	result_output_reg_19,
	result_output_reg_18,
	result_output_reg_17,
	result_output_reg_16,
	result_output_reg_15,
	result_output_reg_14,
	result_output_reg_13,
	result_output_reg_12,
	result_output_reg_11,
	result_output_reg_10,
	result_output_reg_9,
	result_output_reg_8,
	result_output_reg_7,
	result_output_reg_6,
	result_output_reg_5,
	result_output_reg_4,
	result_output_reg_3,
	result_output_reg_2,
	result_output_reg_1,
	result_output_reg_0,
	clock,
	clken)/* synthesis synthesis_greybox=1 */;
input 	[23:0] datab;
input 	[23:0] dataa;
output 	result_output_reg_46;
output 	result_output_reg_23;
output 	result_output_reg_34;
output 	result_output_reg_47;
output 	result_output_reg_24;
output 	result_output_reg_25;
output 	result_output_reg_26;
output 	result_output_reg_27;
output 	result_output_reg_28;
output 	result_output_reg_29;
output 	result_output_reg_30;
output 	result_output_reg_31;
output 	result_output_reg_32;
output 	result_output_reg_33;
output 	result_output_reg_35;
output 	result_output_reg_36;
output 	result_output_reg_37;
output 	result_output_reg_38;
output 	result_output_reg_39;
output 	result_output_reg_40;
output 	result_output_reg_41;
output 	result_output_reg_42;
output 	result_output_reg_43;
output 	result_output_reg_44;
output 	result_output_reg_45;
output 	result_output_reg_22;
output 	result_output_reg_21;
output 	result_output_reg_20;
output 	result_output_reg_19;
output 	result_output_reg_18;
output 	result_output_reg_17;
output 	result_output_reg_16;
output 	result_output_reg_15;
output 	result_output_reg_14;
output 	result_output_reg_13;
output 	result_output_reg_12;
output 	result_output_reg_11;
output 	result_output_reg_10;
output 	result_output_reg_9;
output 	result_output_reg_8;
output 	result_output_reg_7;
output 	result_output_reg_6;
output 	result_output_reg_5;
output 	result_output_reg_4;
output 	result_output_reg_3;
output 	result_output_reg_2;
output 	result_output_reg_1;
output 	result_output_reg_0;
input 	clock;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mult0~8 ;
wire \Mult0~9 ;
wire \Mult0~10 ;
wire \Mult0~11 ;
wire \Mult0~12 ;
wire \Mult0~13 ;
wire \Mult0~14 ;
wire \Mult0~15 ;
wire \Mult0~16 ;
wire \Mult0~17 ;
wire \Mult0~18 ;
wire \Mult0~19 ;
wire \Mult0~20 ;
wire \Mult0~21 ;
wire \Mult0~22 ;
wire \Mult0~23 ;
wire \dataa_input_reg[0]~q ;
wire \dataa_input_reg[1]~q ;
wire \dataa_input_reg[2]~q ;
wire \dataa_input_reg[3]~q ;
wire \dataa_input_reg[4]~q ;
wire \dataa_input_reg[5]~q ;
wire \dataa_input_reg[6]~q ;
wire \dataa_input_reg[7]~q ;
wire \dataa_input_reg[8]~q ;
wire \dataa_input_reg[9]~q ;
wire \dataa_input_reg[10]~q ;
wire \dataa_input_reg[11]~q ;
wire \dataa_input_reg[12]~q ;
wire \dataa_input_reg[13]~q ;
wire \dataa_input_reg[14]~q ;
wire \dataa_input_reg[15]~q ;
wire \dataa_input_reg[16]~q ;
wire \dataa_input_reg[17]~q ;
wire \dataa_input_reg[18]~q ;
wire \dataa_input_reg[19]~q ;
wire \dataa_input_reg[20]~q ;
wire \dataa_input_reg[21]~q ;
wire \dataa_input_reg[22]~q ;
wire \dataa_input_reg[23]~q ;
wire \datab_input_reg[0]~q ;
wire \datab_input_reg[1]~q ;
wire \datab_input_reg[2]~q ;
wire \datab_input_reg[3]~q ;
wire \datab_input_reg[4]~q ;
wire \datab_input_reg[5]~q ;
wire \datab_input_reg[6]~q ;
wire \datab_input_reg[7]~q ;
wire \datab_input_reg[8]~q ;
wire \datab_input_reg[9]~q ;
wire \datab_input_reg[10]~q ;
wire \datab_input_reg[11]~q ;
wire \datab_input_reg[12]~q ;
wire \datab_input_reg[13]~q ;
wire \datab_input_reg[14]~q ;
wire \datab_input_reg[15]~q ;
wire \datab_input_reg[16]~q ;
wire \datab_input_reg[17]~q ;
wire \datab_input_reg[18]~q ;
wire \datab_input_reg[19]~q ;
wire \datab_input_reg[20]~q ;
wire \datab_input_reg[21]~q ;
wire \datab_input_reg[22]~q ;
wire \datab_input_reg[23]~q ;
wire \result_wire[46] ;
wire \result_extra0_reg[46]~q ;
wire \result_wire[23] ;
wire \result_extra0_reg[23]~q ;
wire \result_wire[34] ;
wire \result_extra0_reg[34]~q ;
wire \result_wire[47] ;
wire \result_extra0_reg[47]~q ;
wire \result_wire[24] ;
wire \result_extra0_reg[24]~q ;
wire \result_wire[25] ;
wire \result_extra0_reg[25]~q ;
wire \result_wire[26] ;
wire \result_extra0_reg[26]~q ;
wire \result_wire[27] ;
wire \result_extra0_reg[27]~q ;
wire \result_wire[28] ;
wire \result_extra0_reg[28]~q ;
wire \result_wire[29] ;
wire \result_extra0_reg[29]~q ;
wire \result_wire[30] ;
wire \result_extra0_reg[30]~q ;
wire \result_wire[31] ;
wire \result_extra0_reg[31]~q ;
wire \result_wire[32] ;
wire \result_extra0_reg[32]~q ;
wire \result_wire[33] ;
wire \result_extra0_reg[33]~q ;
wire \result_wire[35] ;
wire \result_extra0_reg[35]~q ;
wire \result_wire[36] ;
wire \result_extra0_reg[36]~q ;
wire \result_wire[37] ;
wire \result_extra0_reg[37]~q ;
wire \result_wire[38] ;
wire \result_extra0_reg[38]~q ;
wire \result_wire[39] ;
wire \result_extra0_reg[39]~q ;
wire \result_wire[40] ;
wire \result_extra0_reg[40]~q ;
wire \result_wire[41] ;
wire \result_extra0_reg[41]~q ;
wire \result_wire[42] ;
wire \result_extra0_reg[42]~q ;
wire \result_wire[43] ;
wire \result_extra0_reg[43]~q ;
wire \result_wire[44] ;
wire \result_extra0_reg[44]~q ;
wire \result_wire[45] ;
wire \result_extra0_reg[45]~q ;
wire \result_wire[22] ;
wire \result_extra0_reg[22]~q ;
wire \result_wire[21] ;
wire \result_extra0_reg[21]~q ;
wire \result_wire[20] ;
wire \result_extra0_reg[20]~q ;
wire \result_wire[19] ;
wire \result_extra0_reg[19]~q ;
wire \result_wire[18] ;
wire \result_extra0_reg[18]~q ;
wire \result_wire[17] ;
wire \result_extra0_reg[17]~q ;
wire \result_wire[16] ;
wire \result_extra0_reg[16]~q ;
wire \result_wire[15] ;
wire \result_extra0_reg[15]~q ;
wire \result_wire[14] ;
wire \result_extra0_reg[14]~q ;
wire \result_wire[13] ;
wire \result_extra0_reg[13]~q ;
wire \result_wire[12] ;
wire \result_extra0_reg[12]~q ;
wire \result_wire[11] ;
wire \result_extra0_reg[11]~q ;
wire \result_wire[10] ;
wire \result_extra0_reg[10]~q ;
wire \result_wire[9] ;
wire \result_extra0_reg[9]~q ;
wire \result_wire[8] ;
wire \result_extra0_reg[8]~q ;
wire \result_wire[7] ;
wire \result_extra0_reg[7]~q ;
wire \result_wire[6] ;
wire \result_extra0_reg[6]~q ;
wire \result_wire[5] ;
wire \result_extra0_reg[5]~q ;
wire \result_wire[4] ;
wire \result_extra0_reg[4]~q ;
wire \result_wire[3] ;
wire \result_extra0_reg[3]~q ;
wire \result_wire[2] ;
wire \result_extra0_reg[2]~q ;
wire \result_wire[1] ;
wire \result_extra0_reg[1]~q ;
wire \result_wire[0] ;
wire \result_extra0_reg[0]~q ;

wire [63:0] \Mult0~mac_RESULTA_bus ;

assign \result_wire[0]  = \Mult0~mac_RESULTA_bus [0];
assign \result_wire[1]  = \Mult0~mac_RESULTA_bus [1];
assign \result_wire[2]  = \Mult0~mac_RESULTA_bus [2];
assign \result_wire[3]  = \Mult0~mac_RESULTA_bus [3];
assign \result_wire[4]  = \Mult0~mac_RESULTA_bus [4];
assign \result_wire[5]  = \Mult0~mac_RESULTA_bus [5];
assign \result_wire[6]  = \Mult0~mac_RESULTA_bus [6];
assign \result_wire[7]  = \Mult0~mac_RESULTA_bus [7];
assign \result_wire[8]  = \Mult0~mac_RESULTA_bus [8];
assign \result_wire[9]  = \Mult0~mac_RESULTA_bus [9];
assign \result_wire[10]  = \Mult0~mac_RESULTA_bus [10];
assign \result_wire[11]  = \Mult0~mac_RESULTA_bus [11];
assign \result_wire[12]  = \Mult0~mac_RESULTA_bus [12];
assign \result_wire[13]  = \Mult0~mac_RESULTA_bus [13];
assign \result_wire[14]  = \Mult0~mac_RESULTA_bus [14];
assign \result_wire[15]  = \Mult0~mac_RESULTA_bus [15];
assign \result_wire[16]  = \Mult0~mac_RESULTA_bus [16];
assign \result_wire[17]  = \Mult0~mac_RESULTA_bus [17];
assign \result_wire[18]  = \Mult0~mac_RESULTA_bus [18];
assign \result_wire[19]  = \Mult0~mac_RESULTA_bus [19];
assign \result_wire[20]  = \Mult0~mac_RESULTA_bus [20];
assign \result_wire[21]  = \Mult0~mac_RESULTA_bus [21];
assign \result_wire[22]  = \Mult0~mac_RESULTA_bus [22];
assign \result_wire[23]  = \Mult0~mac_RESULTA_bus [23];
assign \result_wire[24]  = \Mult0~mac_RESULTA_bus [24];
assign \result_wire[25]  = \Mult0~mac_RESULTA_bus [25];
assign \result_wire[26]  = \Mult0~mac_RESULTA_bus [26];
assign \result_wire[27]  = \Mult0~mac_RESULTA_bus [27];
assign \result_wire[28]  = \Mult0~mac_RESULTA_bus [28];
assign \result_wire[29]  = \Mult0~mac_RESULTA_bus [29];
assign \result_wire[30]  = \Mult0~mac_RESULTA_bus [30];
assign \result_wire[31]  = \Mult0~mac_RESULTA_bus [31];
assign \result_wire[32]  = \Mult0~mac_RESULTA_bus [32];
assign \result_wire[33]  = \Mult0~mac_RESULTA_bus [33];
assign \result_wire[34]  = \Mult0~mac_RESULTA_bus [34];
assign \result_wire[35]  = \Mult0~mac_RESULTA_bus [35];
assign \result_wire[36]  = \Mult0~mac_RESULTA_bus [36];
assign \result_wire[37]  = \Mult0~mac_RESULTA_bus [37];
assign \result_wire[38]  = \Mult0~mac_RESULTA_bus [38];
assign \result_wire[39]  = \Mult0~mac_RESULTA_bus [39];
assign \result_wire[40]  = \Mult0~mac_RESULTA_bus [40];
assign \result_wire[41]  = \Mult0~mac_RESULTA_bus [41];
assign \result_wire[42]  = \Mult0~mac_RESULTA_bus [42];
assign \result_wire[43]  = \Mult0~mac_RESULTA_bus [43];
assign \result_wire[44]  = \Mult0~mac_RESULTA_bus [44];
assign \result_wire[45]  = \Mult0~mac_RESULTA_bus [45];
assign \result_wire[46]  = \Mult0~mac_RESULTA_bus [46];
assign \result_wire[47]  = \Mult0~mac_RESULTA_bus [47];
assign \Mult0~8  = \Mult0~mac_RESULTA_bus [48];
assign \Mult0~9  = \Mult0~mac_RESULTA_bus [49];
assign \Mult0~10  = \Mult0~mac_RESULTA_bus [50];
assign \Mult0~11  = \Mult0~mac_RESULTA_bus [51];
assign \Mult0~12  = \Mult0~mac_RESULTA_bus [52];
assign \Mult0~13  = \Mult0~mac_RESULTA_bus [53];
assign \Mult0~14  = \Mult0~mac_RESULTA_bus [54];
assign \Mult0~15  = \Mult0~mac_RESULTA_bus [55];
assign \Mult0~16  = \Mult0~mac_RESULTA_bus [56];
assign \Mult0~17  = \Mult0~mac_RESULTA_bus [57];
assign \Mult0~18  = \Mult0~mac_RESULTA_bus [58];
assign \Mult0~19  = \Mult0~mac_RESULTA_bus [59];
assign \Mult0~20  = \Mult0~mac_RESULTA_bus [60];
assign \Mult0~21  = \Mult0~mac_RESULTA_bus [61];
assign \Mult0~22  = \Mult0~mac_RESULTA_bus [62];
assign \Mult0~23  = \Mult0~mac_RESULTA_bus [63];

dffeas \result_output_reg[46] (
	.clk(clock),
	.d(\result_extra0_reg[46]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_46),
	.prn(vcc));
defparam \result_output_reg[46] .is_wysiwyg = "true";
defparam \result_output_reg[46] .power_up = "low";

dffeas \result_output_reg[23] (
	.clk(clock),
	.d(\result_extra0_reg[23]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_23),
	.prn(vcc));
defparam \result_output_reg[23] .is_wysiwyg = "true";
defparam \result_output_reg[23] .power_up = "low";

dffeas \result_output_reg[34] (
	.clk(clock),
	.d(\result_extra0_reg[34]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_34),
	.prn(vcc));
defparam \result_output_reg[34] .is_wysiwyg = "true";
defparam \result_output_reg[34] .power_up = "low";

dffeas \result_output_reg[47] (
	.clk(clock),
	.d(\result_extra0_reg[47]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_47),
	.prn(vcc));
defparam \result_output_reg[47] .is_wysiwyg = "true";
defparam \result_output_reg[47] .power_up = "low";

dffeas \result_output_reg[24] (
	.clk(clock),
	.d(\result_extra0_reg[24]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_24),
	.prn(vcc));
defparam \result_output_reg[24] .is_wysiwyg = "true";
defparam \result_output_reg[24] .power_up = "low";

dffeas \result_output_reg[25] (
	.clk(clock),
	.d(\result_extra0_reg[25]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_25),
	.prn(vcc));
defparam \result_output_reg[25] .is_wysiwyg = "true";
defparam \result_output_reg[25] .power_up = "low";

dffeas \result_output_reg[26] (
	.clk(clock),
	.d(\result_extra0_reg[26]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_26),
	.prn(vcc));
defparam \result_output_reg[26] .is_wysiwyg = "true";
defparam \result_output_reg[26] .power_up = "low";

dffeas \result_output_reg[27] (
	.clk(clock),
	.d(\result_extra0_reg[27]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_27),
	.prn(vcc));
defparam \result_output_reg[27] .is_wysiwyg = "true";
defparam \result_output_reg[27] .power_up = "low";

dffeas \result_output_reg[28] (
	.clk(clock),
	.d(\result_extra0_reg[28]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_28),
	.prn(vcc));
defparam \result_output_reg[28] .is_wysiwyg = "true";
defparam \result_output_reg[28] .power_up = "low";

dffeas \result_output_reg[29] (
	.clk(clock),
	.d(\result_extra0_reg[29]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_29),
	.prn(vcc));
defparam \result_output_reg[29] .is_wysiwyg = "true";
defparam \result_output_reg[29] .power_up = "low";

dffeas \result_output_reg[30] (
	.clk(clock),
	.d(\result_extra0_reg[30]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_30),
	.prn(vcc));
defparam \result_output_reg[30] .is_wysiwyg = "true";
defparam \result_output_reg[30] .power_up = "low";

dffeas \result_output_reg[31] (
	.clk(clock),
	.d(\result_extra0_reg[31]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_31),
	.prn(vcc));
defparam \result_output_reg[31] .is_wysiwyg = "true";
defparam \result_output_reg[31] .power_up = "low";

dffeas \result_output_reg[32] (
	.clk(clock),
	.d(\result_extra0_reg[32]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_32),
	.prn(vcc));
defparam \result_output_reg[32] .is_wysiwyg = "true";
defparam \result_output_reg[32] .power_up = "low";

dffeas \result_output_reg[33] (
	.clk(clock),
	.d(\result_extra0_reg[33]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_33),
	.prn(vcc));
defparam \result_output_reg[33] .is_wysiwyg = "true";
defparam \result_output_reg[33] .power_up = "low";

dffeas \result_output_reg[35] (
	.clk(clock),
	.d(\result_extra0_reg[35]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_35),
	.prn(vcc));
defparam \result_output_reg[35] .is_wysiwyg = "true";
defparam \result_output_reg[35] .power_up = "low";

dffeas \result_output_reg[36] (
	.clk(clock),
	.d(\result_extra0_reg[36]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_36),
	.prn(vcc));
defparam \result_output_reg[36] .is_wysiwyg = "true";
defparam \result_output_reg[36] .power_up = "low";

dffeas \result_output_reg[37] (
	.clk(clock),
	.d(\result_extra0_reg[37]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_37),
	.prn(vcc));
defparam \result_output_reg[37] .is_wysiwyg = "true";
defparam \result_output_reg[37] .power_up = "low";

dffeas \result_output_reg[38] (
	.clk(clock),
	.d(\result_extra0_reg[38]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_38),
	.prn(vcc));
defparam \result_output_reg[38] .is_wysiwyg = "true";
defparam \result_output_reg[38] .power_up = "low";

dffeas \result_output_reg[39] (
	.clk(clock),
	.d(\result_extra0_reg[39]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_39),
	.prn(vcc));
defparam \result_output_reg[39] .is_wysiwyg = "true";
defparam \result_output_reg[39] .power_up = "low";

dffeas \result_output_reg[40] (
	.clk(clock),
	.d(\result_extra0_reg[40]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_40),
	.prn(vcc));
defparam \result_output_reg[40] .is_wysiwyg = "true";
defparam \result_output_reg[40] .power_up = "low";

dffeas \result_output_reg[41] (
	.clk(clock),
	.d(\result_extra0_reg[41]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_41),
	.prn(vcc));
defparam \result_output_reg[41] .is_wysiwyg = "true";
defparam \result_output_reg[41] .power_up = "low";

dffeas \result_output_reg[42] (
	.clk(clock),
	.d(\result_extra0_reg[42]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_42),
	.prn(vcc));
defparam \result_output_reg[42] .is_wysiwyg = "true";
defparam \result_output_reg[42] .power_up = "low";

dffeas \result_output_reg[43] (
	.clk(clock),
	.d(\result_extra0_reg[43]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_43),
	.prn(vcc));
defparam \result_output_reg[43] .is_wysiwyg = "true";
defparam \result_output_reg[43] .power_up = "low";

dffeas \result_output_reg[44] (
	.clk(clock),
	.d(\result_extra0_reg[44]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_44),
	.prn(vcc));
defparam \result_output_reg[44] .is_wysiwyg = "true";
defparam \result_output_reg[44] .power_up = "low";

dffeas \result_output_reg[45] (
	.clk(clock),
	.d(\result_extra0_reg[45]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_45),
	.prn(vcc));
defparam \result_output_reg[45] .is_wysiwyg = "true";
defparam \result_output_reg[45] .power_up = "low";

dffeas \result_output_reg[22] (
	.clk(clock),
	.d(\result_extra0_reg[22]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_22),
	.prn(vcc));
defparam \result_output_reg[22] .is_wysiwyg = "true";
defparam \result_output_reg[22] .power_up = "low";

dffeas \result_output_reg[21] (
	.clk(clock),
	.d(\result_extra0_reg[21]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_21),
	.prn(vcc));
defparam \result_output_reg[21] .is_wysiwyg = "true";
defparam \result_output_reg[21] .power_up = "low";

dffeas \result_output_reg[20] (
	.clk(clock),
	.d(\result_extra0_reg[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_20),
	.prn(vcc));
defparam \result_output_reg[20] .is_wysiwyg = "true";
defparam \result_output_reg[20] .power_up = "low";

dffeas \result_output_reg[19] (
	.clk(clock),
	.d(\result_extra0_reg[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_19),
	.prn(vcc));
defparam \result_output_reg[19] .is_wysiwyg = "true";
defparam \result_output_reg[19] .power_up = "low";

dffeas \result_output_reg[18] (
	.clk(clock),
	.d(\result_extra0_reg[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_18),
	.prn(vcc));
defparam \result_output_reg[18] .is_wysiwyg = "true";
defparam \result_output_reg[18] .power_up = "low";

dffeas \result_output_reg[17] (
	.clk(clock),
	.d(\result_extra0_reg[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_17),
	.prn(vcc));
defparam \result_output_reg[17] .is_wysiwyg = "true";
defparam \result_output_reg[17] .power_up = "low";

dffeas \result_output_reg[16] (
	.clk(clock),
	.d(\result_extra0_reg[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_16),
	.prn(vcc));
defparam \result_output_reg[16] .is_wysiwyg = "true";
defparam \result_output_reg[16] .power_up = "low";

dffeas \result_output_reg[15] (
	.clk(clock),
	.d(\result_extra0_reg[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_15),
	.prn(vcc));
defparam \result_output_reg[15] .is_wysiwyg = "true";
defparam \result_output_reg[15] .power_up = "low";

dffeas \result_output_reg[14] (
	.clk(clock),
	.d(\result_extra0_reg[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_14),
	.prn(vcc));
defparam \result_output_reg[14] .is_wysiwyg = "true";
defparam \result_output_reg[14] .power_up = "low";

dffeas \result_output_reg[13] (
	.clk(clock),
	.d(\result_extra0_reg[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_13),
	.prn(vcc));
defparam \result_output_reg[13] .is_wysiwyg = "true";
defparam \result_output_reg[13] .power_up = "low";

dffeas \result_output_reg[12] (
	.clk(clock),
	.d(\result_extra0_reg[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_12),
	.prn(vcc));
defparam \result_output_reg[12] .is_wysiwyg = "true";
defparam \result_output_reg[12] .power_up = "low";

dffeas \result_output_reg[11] (
	.clk(clock),
	.d(\result_extra0_reg[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_11),
	.prn(vcc));
defparam \result_output_reg[11] .is_wysiwyg = "true";
defparam \result_output_reg[11] .power_up = "low";

dffeas \result_output_reg[10] (
	.clk(clock),
	.d(\result_extra0_reg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_10),
	.prn(vcc));
defparam \result_output_reg[10] .is_wysiwyg = "true";
defparam \result_output_reg[10] .power_up = "low";

dffeas \result_output_reg[9] (
	.clk(clock),
	.d(\result_extra0_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_9),
	.prn(vcc));
defparam \result_output_reg[9] .is_wysiwyg = "true";
defparam \result_output_reg[9] .power_up = "low";

dffeas \result_output_reg[8] (
	.clk(clock),
	.d(\result_extra0_reg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_8),
	.prn(vcc));
defparam \result_output_reg[8] .is_wysiwyg = "true";
defparam \result_output_reg[8] .power_up = "low";

dffeas \result_output_reg[7] (
	.clk(clock),
	.d(\result_extra0_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_7),
	.prn(vcc));
defparam \result_output_reg[7] .is_wysiwyg = "true";
defparam \result_output_reg[7] .power_up = "low";

dffeas \result_output_reg[6] (
	.clk(clock),
	.d(\result_extra0_reg[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_6),
	.prn(vcc));
defparam \result_output_reg[6] .is_wysiwyg = "true";
defparam \result_output_reg[6] .power_up = "low";

dffeas \result_output_reg[5] (
	.clk(clock),
	.d(\result_extra0_reg[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_5),
	.prn(vcc));
defparam \result_output_reg[5] .is_wysiwyg = "true";
defparam \result_output_reg[5] .power_up = "low";

dffeas \result_output_reg[4] (
	.clk(clock),
	.d(\result_extra0_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_4),
	.prn(vcc));
defparam \result_output_reg[4] .is_wysiwyg = "true";
defparam \result_output_reg[4] .power_up = "low";

dffeas \result_output_reg[3] (
	.clk(clock),
	.d(\result_extra0_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_3),
	.prn(vcc));
defparam \result_output_reg[3] .is_wysiwyg = "true";
defparam \result_output_reg[3] .power_up = "low";

dffeas \result_output_reg[2] (
	.clk(clock),
	.d(\result_extra0_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_2),
	.prn(vcc));
defparam \result_output_reg[2] .is_wysiwyg = "true";
defparam \result_output_reg[2] .power_up = "low";

dffeas \result_output_reg[1] (
	.clk(clock),
	.d(\result_extra0_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_1),
	.prn(vcc));
defparam \result_output_reg[1] .is_wysiwyg = "true";
defparam \result_output_reg[1] .power_up = "low";

dffeas \result_output_reg[0] (
	.clk(clock),
	.d(\result_extra0_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(result_output_reg_0),
	.prn(vcc));
defparam \result_output_reg[0] .is_wysiwyg = "true";
defparam \result_output_reg[0] .power_up = "low";

dffeas \dataa_input_reg[0] (
	.clk(clock),
	.d(dataa[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[0]~q ),
	.prn(vcc));
defparam \dataa_input_reg[0] .is_wysiwyg = "true";
defparam \dataa_input_reg[0] .power_up = "low";

dffeas \dataa_input_reg[1] (
	.clk(clock),
	.d(dataa[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[1]~q ),
	.prn(vcc));
defparam \dataa_input_reg[1] .is_wysiwyg = "true";
defparam \dataa_input_reg[1] .power_up = "low";

dffeas \dataa_input_reg[2] (
	.clk(clock),
	.d(dataa[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[2]~q ),
	.prn(vcc));
defparam \dataa_input_reg[2] .is_wysiwyg = "true";
defparam \dataa_input_reg[2] .power_up = "low";

dffeas \dataa_input_reg[3] (
	.clk(clock),
	.d(dataa[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[3]~q ),
	.prn(vcc));
defparam \dataa_input_reg[3] .is_wysiwyg = "true";
defparam \dataa_input_reg[3] .power_up = "low";

dffeas \dataa_input_reg[4] (
	.clk(clock),
	.d(dataa[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[4]~q ),
	.prn(vcc));
defparam \dataa_input_reg[4] .is_wysiwyg = "true";
defparam \dataa_input_reg[4] .power_up = "low";

dffeas \dataa_input_reg[5] (
	.clk(clock),
	.d(dataa[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[5]~q ),
	.prn(vcc));
defparam \dataa_input_reg[5] .is_wysiwyg = "true";
defparam \dataa_input_reg[5] .power_up = "low";

dffeas \dataa_input_reg[6] (
	.clk(clock),
	.d(dataa[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[6]~q ),
	.prn(vcc));
defparam \dataa_input_reg[6] .is_wysiwyg = "true";
defparam \dataa_input_reg[6] .power_up = "low";

dffeas \dataa_input_reg[7] (
	.clk(clock),
	.d(dataa[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[7]~q ),
	.prn(vcc));
defparam \dataa_input_reg[7] .is_wysiwyg = "true";
defparam \dataa_input_reg[7] .power_up = "low";

dffeas \dataa_input_reg[8] (
	.clk(clock),
	.d(dataa[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[8]~q ),
	.prn(vcc));
defparam \dataa_input_reg[8] .is_wysiwyg = "true";
defparam \dataa_input_reg[8] .power_up = "low";

dffeas \dataa_input_reg[9] (
	.clk(clock),
	.d(dataa[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[9]~q ),
	.prn(vcc));
defparam \dataa_input_reg[9] .is_wysiwyg = "true";
defparam \dataa_input_reg[9] .power_up = "low";

dffeas \dataa_input_reg[10] (
	.clk(clock),
	.d(dataa[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[10]~q ),
	.prn(vcc));
defparam \dataa_input_reg[10] .is_wysiwyg = "true";
defparam \dataa_input_reg[10] .power_up = "low";

dffeas \dataa_input_reg[11] (
	.clk(clock),
	.d(dataa[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[11]~q ),
	.prn(vcc));
defparam \dataa_input_reg[11] .is_wysiwyg = "true";
defparam \dataa_input_reg[11] .power_up = "low";

dffeas \dataa_input_reg[12] (
	.clk(clock),
	.d(dataa[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[12]~q ),
	.prn(vcc));
defparam \dataa_input_reg[12] .is_wysiwyg = "true";
defparam \dataa_input_reg[12] .power_up = "low";

dffeas \dataa_input_reg[13] (
	.clk(clock),
	.d(dataa[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[13]~q ),
	.prn(vcc));
defparam \dataa_input_reg[13] .is_wysiwyg = "true";
defparam \dataa_input_reg[13] .power_up = "low";

dffeas \dataa_input_reg[14] (
	.clk(clock),
	.d(dataa[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[14]~q ),
	.prn(vcc));
defparam \dataa_input_reg[14] .is_wysiwyg = "true";
defparam \dataa_input_reg[14] .power_up = "low";

dffeas \dataa_input_reg[15] (
	.clk(clock),
	.d(dataa[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[15]~q ),
	.prn(vcc));
defparam \dataa_input_reg[15] .is_wysiwyg = "true";
defparam \dataa_input_reg[15] .power_up = "low";

dffeas \dataa_input_reg[16] (
	.clk(clock),
	.d(dataa[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[16]~q ),
	.prn(vcc));
defparam \dataa_input_reg[16] .is_wysiwyg = "true";
defparam \dataa_input_reg[16] .power_up = "low";

dffeas \dataa_input_reg[17] (
	.clk(clock),
	.d(dataa[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[17]~q ),
	.prn(vcc));
defparam \dataa_input_reg[17] .is_wysiwyg = "true";
defparam \dataa_input_reg[17] .power_up = "low";

dffeas \dataa_input_reg[18] (
	.clk(clock),
	.d(dataa[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[18]~q ),
	.prn(vcc));
defparam \dataa_input_reg[18] .is_wysiwyg = "true";
defparam \dataa_input_reg[18] .power_up = "low";

dffeas \dataa_input_reg[19] (
	.clk(clock),
	.d(dataa[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[19]~q ),
	.prn(vcc));
defparam \dataa_input_reg[19] .is_wysiwyg = "true";
defparam \dataa_input_reg[19] .power_up = "low";

dffeas \dataa_input_reg[20] (
	.clk(clock),
	.d(dataa[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[20]~q ),
	.prn(vcc));
defparam \dataa_input_reg[20] .is_wysiwyg = "true";
defparam \dataa_input_reg[20] .power_up = "low";

dffeas \dataa_input_reg[21] (
	.clk(clock),
	.d(dataa[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[21]~q ),
	.prn(vcc));
defparam \dataa_input_reg[21] .is_wysiwyg = "true";
defparam \dataa_input_reg[21] .power_up = "low";

dffeas \dataa_input_reg[22] (
	.clk(clock),
	.d(dataa[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[22]~q ),
	.prn(vcc));
defparam \dataa_input_reg[22] .is_wysiwyg = "true";
defparam \dataa_input_reg[22] .power_up = "low";

dffeas \dataa_input_reg[23] (
	.clk(clock),
	.d(dataa[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dataa_input_reg[23]~q ),
	.prn(vcc));
defparam \dataa_input_reg[23] .is_wysiwyg = "true";
defparam \dataa_input_reg[23] .power_up = "low";

dffeas \datab_input_reg[0] (
	.clk(clock),
	.d(datab[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[0]~q ),
	.prn(vcc));
defparam \datab_input_reg[0] .is_wysiwyg = "true";
defparam \datab_input_reg[0] .power_up = "low";

dffeas \datab_input_reg[1] (
	.clk(clock),
	.d(datab[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[1]~q ),
	.prn(vcc));
defparam \datab_input_reg[1] .is_wysiwyg = "true";
defparam \datab_input_reg[1] .power_up = "low";

dffeas \datab_input_reg[2] (
	.clk(clock),
	.d(datab[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[2]~q ),
	.prn(vcc));
defparam \datab_input_reg[2] .is_wysiwyg = "true";
defparam \datab_input_reg[2] .power_up = "low";

dffeas \datab_input_reg[3] (
	.clk(clock),
	.d(datab[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[3]~q ),
	.prn(vcc));
defparam \datab_input_reg[3] .is_wysiwyg = "true";
defparam \datab_input_reg[3] .power_up = "low";

dffeas \datab_input_reg[4] (
	.clk(clock),
	.d(datab[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[4]~q ),
	.prn(vcc));
defparam \datab_input_reg[4] .is_wysiwyg = "true";
defparam \datab_input_reg[4] .power_up = "low";

dffeas \datab_input_reg[5] (
	.clk(clock),
	.d(datab[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[5]~q ),
	.prn(vcc));
defparam \datab_input_reg[5] .is_wysiwyg = "true";
defparam \datab_input_reg[5] .power_up = "low";

dffeas \datab_input_reg[6] (
	.clk(clock),
	.d(datab[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[6]~q ),
	.prn(vcc));
defparam \datab_input_reg[6] .is_wysiwyg = "true";
defparam \datab_input_reg[6] .power_up = "low";

dffeas \datab_input_reg[7] (
	.clk(clock),
	.d(datab[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[7]~q ),
	.prn(vcc));
defparam \datab_input_reg[7] .is_wysiwyg = "true";
defparam \datab_input_reg[7] .power_up = "low";

dffeas \datab_input_reg[8] (
	.clk(clock),
	.d(datab[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[8]~q ),
	.prn(vcc));
defparam \datab_input_reg[8] .is_wysiwyg = "true";
defparam \datab_input_reg[8] .power_up = "low";

dffeas \datab_input_reg[9] (
	.clk(clock),
	.d(datab[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[9]~q ),
	.prn(vcc));
defparam \datab_input_reg[9] .is_wysiwyg = "true";
defparam \datab_input_reg[9] .power_up = "low";

dffeas \datab_input_reg[10] (
	.clk(clock),
	.d(datab[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[10]~q ),
	.prn(vcc));
defparam \datab_input_reg[10] .is_wysiwyg = "true";
defparam \datab_input_reg[10] .power_up = "low";

dffeas \datab_input_reg[11] (
	.clk(clock),
	.d(datab[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[11]~q ),
	.prn(vcc));
defparam \datab_input_reg[11] .is_wysiwyg = "true";
defparam \datab_input_reg[11] .power_up = "low";

dffeas \datab_input_reg[12] (
	.clk(clock),
	.d(datab[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[12]~q ),
	.prn(vcc));
defparam \datab_input_reg[12] .is_wysiwyg = "true";
defparam \datab_input_reg[12] .power_up = "low";

dffeas \datab_input_reg[13] (
	.clk(clock),
	.d(datab[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[13]~q ),
	.prn(vcc));
defparam \datab_input_reg[13] .is_wysiwyg = "true";
defparam \datab_input_reg[13] .power_up = "low";

dffeas \datab_input_reg[14] (
	.clk(clock),
	.d(datab[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[14]~q ),
	.prn(vcc));
defparam \datab_input_reg[14] .is_wysiwyg = "true";
defparam \datab_input_reg[14] .power_up = "low";

dffeas \datab_input_reg[15] (
	.clk(clock),
	.d(datab[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[15]~q ),
	.prn(vcc));
defparam \datab_input_reg[15] .is_wysiwyg = "true";
defparam \datab_input_reg[15] .power_up = "low";

dffeas \datab_input_reg[16] (
	.clk(clock),
	.d(datab[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[16]~q ),
	.prn(vcc));
defparam \datab_input_reg[16] .is_wysiwyg = "true";
defparam \datab_input_reg[16] .power_up = "low";

dffeas \datab_input_reg[17] (
	.clk(clock),
	.d(datab[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[17]~q ),
	.prn(vcc));
defparam \datab_input_reg[17] .is_wysiwyg = "true";
defparam \datab_input_reg[17] .power_up = "low";

dffeas \datab_input_reg[18] (
	.clk(clock),
	.d(datab[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[18]~q ),
	.prn(vcc));
defparam \datab_input_reg[18] .is_wysiwyg = "true";
defparam \datab_input_reg[18] .power_up = "low";

dffeas \datab_input_reg[19] (
	.clk(clock),
	.d(datab[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[19]~q ),
	.prn(vcc));
defparam \datab_input_reg[19] .is_wysiwyg = "true";
defparam \datab_input_reg[19] .power_up = "low";

dffeas \datab_input_reg[20] (
	.clk(clock),
	.d(datab[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[20]~q ),
	.prn(vcc));
defparam \datab_input_reg[20] .is_wysiwyg = "true";
defparam \datab_input_reg[20] .power_up = "low";

dffeas \datab_input_reg[21] (
	.clk(clock),
	.d(datab[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[21]~q ),
	.prn(vcc));
defparam \datab_input_reg[21] .is_wysiwyg = "true";
defparam \datab_input_reg[21] .power_up = "low";

dffeas \datab_input_reg[22] (
	.clk(clock),
	.d(datab[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[22]~q ),
	.prn(vcc));
defparam \datab_input_reg[22] .is_wysiwyg = "true";
defparam \datab_input_reg[22] .power_up = "low";

dffeas \datab_input_reg[23] (
	.clk(clock),
	.d(datab[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\datab_input_reg[23]~q ),
	.prn(vcc));
defparam \datab_input_reg[23] .is_wysiwyg = "true";
defparam \datab_input_reg[23] .power_up = "low";

cyclonev_mac \Mult0~mac (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,\dataa_input_reg[23]~q ,\dataa_input_reg[22]~q ,\dataa_input_reg[21]~q ,\dataa_input_reg[20]~q ,\dataa_input_reg[19]~q ,\dataa_input_reg[18]~q ,\dataa_input_reg[17]~q ,\dataa_input_reg[16]~q ,\dataa_input_reg[15]~q ,\dataa_input_reg[14]~q ,
\dataa_input_reg[13]~q ,\dataa_input_reg[12]~q ,\dataa_input_reg[11]~q ,\dataa_input_reg[10]~q ,\dataa_input_reg[9]~q ,\dataa_input_reg[8]~q ,\dataa_input_reg[7]~q ,\dataa_input_reg[6]~q ,\dataa_input_reg[5]~q ,\dataa_input_reg[4]~q ,\dataa_input_reg[3]~q ,
\dataa_input_reg[2]~q ,\dataa_input_reg[1]~q ,\dataa_input_reg[0]~q }),
	.ay({gnd,gnd,gnd,\datab_input_reg[23]~q ,\datab_input_reg[22]~q ,\datab_input_reg[21]~q ,\datab_input_reg[20]~q ,\datab_input_reg[19]~q ,\datab_input_reg[18]~q ,\datab_input_reg[17]~q ,\datab_input_reg[16]~q ,\datab_input_reg[15]~q ,\datab_input_reg[14]~q ,
\datab_input_reg[13]~q ,\datab_input_reg[12]~q ,\datab_input_reg[11]~q ,\datab_input_reg[10]~q ,\datab_input_reg[9]~q ,\datab_input_reg[8]~q ,\datab_input_reg[7]~q ,\datab_input_reg[6]~q ,\datab_input_reg[5]~q ,\datab_input_reg[4]~q ,\datab_input_reg[3]~q ,
\datab_input_reg[2]~q ,\datab_input_reg[1]~q ,\datab_input_reg[0]~q }),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Mult0~mac_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Mult0~mac .accumulate_clock = "none";
defparam \Mult0~mac .ax_clock = "none";
defparam \Mult0~mac .ax_width = 24;
defparam \Mult0~mac .ay_scan_in_clock = "none";
defparam \Mult0~mac .ay_scan_in_width = 24;
defparam \Mult0~mac .ay_use_scan_in = "false";
defparam \Mult0~mac .az_clock = "none";
defparam \Mult0~mac .bx_clock = "none";
defparam \Mult0~mac .by_clock = "none";
defparam \Mult0~mac .by_use_scan_in = "false";
defparam \Mult0~mac .bz_clock = "none";
defparam \Mult0~mac .coef_a_0 = 0;
defparam \Mult0~mac .coef_a_1 = 0;
defparam \Mult0~mac .coef_a_2 = 0;
defparam \Mult0~mac .coef_a_3 = 0;
defparam \Mult0~mac .coef_a_4 = 0;
defparam \Mult0~mac .coef_a_5 = 0;
defparam \Mult0~mac .coef_a_6 = 0;
defparam \Mult0~mac .coef_a_7 = 0;
defparam \Mult0~mac .coef_b_0 = 0;
defparam \Mult0~mac .coef_b_1 = 0;
defparam \Mult0~mac .coef_b_2 = 0;
defparam \Mult0~mac .coef_b_3 = 0;
defparam \Mult0~mac .coef_b_4 = 0;
defparam \Mult0~mac .coef_b_5 = 0;
defparam \Mult0~mac .coef_b_6 = 0;
defparam \Mult0~mac .coef_b_7 = 0;
defparam \Mult0~mac .coef_sel_a_clock = "none";
defparam \Mult0~mac .coef_sel_b_clock = "none";
defparam \Mult0~mac .delay_scan_out_ay = "false";
defparam \Mult0~mac .delay_scan_out_by = "false";
defparam \Mult0~mac .enable_double_accum = "false";
defparam \Mult0~mac .load_const_clock = "none";
defparam \Mult0~mac .load_const_value = 0;
defparam \Mult0~mac .mode_sub_location = 0;
defparam \Mult0~mac .negate_clock = "none";
defparam \Mult0~mac .operand_source_max = "input";
defparam \Mult0~mac .operand_source_may = "input";
defparam \Mult0~mac .operand_source_mbx = "input";
defparam \Mult0~mac .operand_source_mby = "input";
defparam \Mult0~mac .operation_mode = "m27x27";
defparam \Mult0~mac .output_clock = "none";
defparam \Mult0~mac .preadder_subtract_a = "false";
defparam \Mult0~mac .preadder_subtract_b = "false";
defparam \Mult0~mac .result_a_width = 64;
defparam \Mult0~mac .signed_max = "true";
defparam \Mult0~mac .signed_may = "true";
defparam \Mult0~mac .signed_mbx = "false";
defparam \Mult0~mac .signed_mby = "false";
defparam \Mult0~mac .sub_clock = "none";
defparam \Mult0~mac .use_chainadder = "false";

dffeas \result_extra0_reg[46] (
	.clk(clock),
	.d(\result_wire[46] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[46]~q ),
	.prn(vcc));
defparam \result_extra0_reg[46] .is_wysiwyg = "true";
defparam \result_extra0_reg[46] .power_up = "low";

dffeas \result_extra0_reg[23] (
	.clk(clock),
	.d(\result_wire[23] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[23]~q ),
	.prn(vcc));
defparam \result_extra0_reg[23] .is_wysiwyg = "true";
defparam \result_extra0_reg[23] .power_up = "low";

dffeas \result_extra0_reg[34] (
	.clk(clock),
	.d(\result_wire[34] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[34]~q ),
	.prn(vcc));
defparam \result_extra0_reg[34] .is_wysiwyg = "true";
defparam \result_extra0_reg[34] .power_up = "low";

dffeas \result_extra0_reg[47] (
	.clk(clock),
	.d(\result_wire[47] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[47]~q ),
	.prn(vcc));
defparam \result_extra0_reg[47] .is_wysiwyg = "true";
defparam \result_extra0_reg[47] .power_up = "low";

dffeas \result_extra0_reg[24] (
	.clk(clock),
	.d(\result_wire[24] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[24]~q ),
	.prn(vcc));
defparam \result_extra0_reg[24] .is_wysiwyg = "true";
defparam \result_extra0_reg[24] .power_up = "low";

dffeas \result_extra0_reg[25] (
	.clk(clock),
	.d(\result_wire[25] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[25]~q ),
	.prn(vcc));
defparam \result_extra0_reg[25] .is_wysiwyg = "true";
defparam \result_extra0_reg[25] .power_up = "low";

dffeas \result_extra0_reg[26] (
	.clk(clock),
	.d(\result_wire[26] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[26]~q ),
	.prn(vcc));
defparam \result_extra0_reg[26] .is_wysiwyg = "true";
defparam \result_extra0_reg[26] .power_up = "low";

dffeas \result_extra0_reg[27] (
	.clk(clock),
	.d(\result_wire[27] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[27]~q ),
	.prn(vcc));
defparam \result_extra0_reg[27] .is_wysiwyg = "true";
defparam \result_extra0_reg[27] .power_up = "low";

dffeas \result_extra0_reg[28] (
	.clk(clock),
	.d(\result_wire[28] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[28]~q ),
	.prn(vcc));
defparam \result_extra0_reg[28] .is_wysiwyg = "true";
defparam \result_extra0_reg[28] .power_up = "low";

dffeas \result_extra0_reg[29] (
	.clk(clock),
	.d(\result_wire[29] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[29]~q ),
	.prn(vcc));
defparam \result_extra0_reg[29] .is_wysiwyg = "true";
defparam \result_extra0_reg[29] .power_up = "low";

dffeas \result_extra0_reg[30] (
	.clk(clock),
	.d(\result_wire[30] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[30]~q ),
	.prn(vcc));
defparam \result_extra0_reg[30] .is_wysiwyg = "true";
defparam \result_extra0_reg[30] .power_up = "low";

dffeas \result_extra0_reg[31] (
	.clk(clock),
	.d(\result_wire[31] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[31]~q ),
	.prn(vcc));
defparam \result_extra0_reg[31] .is_wysiwyg = "true";
defparam \result_extra0_reg[31] .power_up = "low";

dffeas \result_extra0_reg[32] (
	.clk(clock),
	.d(\result_wire[32] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[32]~q ),
	.prn(vcc));
defparam \result_extra0_reg[32] .is_wysiwyg = "true";
defparam \result_extra0_reg[32] .power_up = "low";

dffeas \result_extra0_reg[33] (
	.clk(clock),
	.d(\result_wire[33] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[33]~q ),
	.prn(vcc));
defparam \result_extra0_reg[33] .is_wysiwyg = "true";
defparam \result_extra0_reg[33] .power_up = "low";

dffeas \result_extra0_reg[35] (
	.clk(clock),
	.d(\result_wire[35] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[35]~q ),
	.prn(vcc));
defparam \result_extra0_reg[35] .is_wysiwyg = "true";
defparam \result_extra0_reg[35] .power_up = "low";

dffeas \result_extra0_reg[36] (
	.clk(clock),
	.d(\result_wire[36] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[36]~q ),
	.prn(vcc));
defparam \result_extra0_reg[36] .is_wysiwyg = "true";
defparam \result_extra0_reg[36] .power_up = "low";

dffeas \result_extra0_reg[37] (
	.clk(clock),
	.d(\result_wire[37] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[37]~q ),
	.prn(vcc));
defparam \result_extra0_reg[37] .is_wysiwyg = "true";
defparam \result_extra0_reg[37] .power_up = "low";

dffeas \result_extra0_reg[38] (
	.clk(clock),
	.d(\result_wire[38] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[38]~q ),
	.prn(vcc));
defparam \result_extra0_reg[38] .is_wysiwyg = "true";
defparam \result_extra0_reg[38] .power_up = "low";

dffeas \result_extra0_reg[39] (
	.clk(clock),
	.d(\result_wire[39] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[39]~q ),
	.prn(vcc));
defparam \result_extra0_reg[39] .is_wysiwyg = "true";
defparam \result_extra0_reg[39] .power_up = "low";

dffeas \result_extra0_reg[40] (
	.clk(clock),
	.d(\result_wire[40] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[40]~q ),
	.prn(vcc));
defparam \result_extra0_reg[40] .is_wysiwyg = "true";
defparam \result_extra0_reg[40] .power_up = "low";

dffeas \result_extra0_reg[41] (
	.clk(clock),
	.d(\result_wire[41] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[41]~q ),
	.prn(vcc));
defparam \result_extra0_reg[41] .is_wysiwyg = "true";
defparam \result_extra0_reg[41] .power_up = "low";

dffeas \result_extra0_reg[42] (
	.clk(clock),
	.d(\result_wire[42] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[42]~q ),
	.prn(vcc));
defparam \result_extra0_reg[42] .is_wysiwyg = "true";
defparam \result_extra0_reg[42] .power_up = "low";

dffeas \result_extra0_reg[43] (
	.clk(clock),
	.d(\result_wire[43] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[43]~q ),
	.prn(vcc));
defparam \result_extra0_reg[43] .is_wysiwyg = "true";
defparam \result_extra0_reg[43] .power_up = "low";

dffeas \result_extra0_reg[44] (
	.clk(clock),
	.d(\result_wire[44] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[44]~q ),
	.prn(vcc));
defparam \result_extra0_reg[44] .is_wysiwyg = "true";
defparam \result_extra0_reg[44] .power_up = "low";

dffeas \result_extra0_reg[45] (
	.clk(clock),
	.d(\result_wire[45] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[45]~q ),
	.prn(vcc));
defparam \result_extra0_reg[45] .is_wysiwyg = "true";
defparam \result_extra0_reg[45] .power_up = "low";

dffeas \result_extra0_reg[22] (
	.clk(clock),
	.d(\result_wire[22] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[22]~q ),
	.prn(vcc));
defparam \result_extra0_reg[22] .is_wysiwyg = "true";
defparam \result_extra0_reg[22] .power_up = "low";

dffeas \result_extra0_reg[21] (
	.clk(clock),
	.d(\result_wire[21] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[21]~q ),
	.prn(vcc));
defparam \result_extra0_reg[21] .is_wysiwyg = "true";
defparam \result_extra0_reg[21] .power_up = "low";

dffeas \result_extra0_reg[20] (
	.clk(clock),
	.d(\result_wire[20] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[20]~q ),
	.prn(vcc));
defparam \result_extra0_reg[20] .is_wysiwyg = "true";
defparam \result_extra0_reg[20] .power_up = "low";

dffeas \result_extra0_reg[19] (
	.clk(clock),
	.d(\result_wire[19] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[19]~q ),
	.prn(vcc));
defparam \result_extra0_reg[19] .is_wysiwyg = "true";
defparam \result_extra0_reg[19] .power_up = "low";

dffeas \result_extra0_reg[18] (
	.clk(clock),
	.d(\result_wire[18] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[18]~q ),
	.prn(vcc));
defparam \result_extra0_reg[18] .is_wysiwyg = "true";
defparam \result_extra0_reg[18] .power_up = "low";

dffeas \result_extra0_reg[17] (
	.clk(clock),
	.d(\result_wire[17] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[17]~q ),
	.prn(vcc));
defparam \result_extra0_reg[17] .is_wysiwyg = "true";
defparam \result_extra0_reg[17] .power_up = "low";

dffeas \result_extra0_reg[16] (
	.clk(clock),
	.d(\result_wire[16] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[16]~q ),
	.prn(vcc));
defparam \result_extra0_reg[16] .is_wysiwyg = "true";
defparam \result_extra0_reg[16] .power_up = "low";

dffeas \result_extra0_reg[15] (
	.clk(clock),
	.d(\result_wire[15] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[15]~q ),
	.prn(vcc));
defparam \result_extra0_reg[15] .is_wysiwyg = "true";
defparam \result_extra0_reg[15] .power_up = "low";

dffeas \result_extra0_reg[14] (
	.clk(clock),
	.d(\result_wire[14] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[14]~q ),
	.prn(vcc));
defparam \result_extra0_reg[14] .is_wysiwyg = "true";
defparam \result_extra0_reg[14] .power_up = "low";

dffeas \result_extra0_reg[13] (
	.clk(clock),
	.d(\result_wire[13] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[13]~q ),
	.prn(vcc));
defparam \result_extra0_reg[13] .is_wysiwyg = "true";
defparam \result_extra0_reg[13] .power_up = "low";

dffeas \result_extra0_reg[12] (
	.clk(clock),
	.d(\result_wire[12] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[12]~q ),
	.prn(vcc));
defparam \result_extra0_reg[12] .is_wysiwyg = "true";
defparam \result_extra0_reg[12] .power_up = "low";

dffeas \result_extra0_reg[11] (
	.clk(clock),
	.d(\result_wire[11] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[11]~q ),
	.prn(vcc));
defparam \result_extra0_reg[11] .is_wysiwyg = "true";
defparam \result_extra0_reg[11] .power_up = "low";

dffeas \result_extra0_reg[10] (
	.clk(clock),
	.d(\result_wire[10] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[10]~q ),
	.prn(vcc));
defparam \result_extra0_reg[10] .is_wysiwyg = "true";
defparam \result_extra0_reg[10] .power_up = "low";

dffeas \result_extra0_reg[9] (
	.clk(clock),
	.d(\result_wire[9] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[9]~q ),
	.prn(vcc));
defparam \result_extra0_reg[9] .is_wysiwyg = "true";
defparam \result_extra0_reg[9] .power_up = "low";

dffeas \result_extra0_reg[8] (
	.clk(clock),
	.d(\result_wire[8] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[8]~q ),
	.prn(vcc));
defparam \result_extra0_reg[8] .is_wysiwyg = "true";
defparam \result_extra0_reg[8] .power_up = "low";

dffeas \result_extra0_reg[7] (
	.clk(clock),
	.d(\result_wire[7] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[7]~q ),
	.prn(vcc));
defparam \result_extra0_reg[7] .is_wysiwyg = "true";
defparam \result_extra0_reg[7] .power_up = "low";

dffeas \result_extra0_reg[6] (
	.clk(clock),
	.d(\result_wire[6] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[6]~q ),
	.prn(vcc));
defparam \result_extra0_reg[6] .is_wysiwyg = "true";
defparam \result_extra0_reg[6] .power_up = "low";

dffeas \result_extra0_reg[5] (
	.clk(clock),
	.d(\result_wire[5] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[5]~q ),
	.prn(vcc));
defparam \result_extra0_reg[5] .is_wysiwyg = "true";
defparam \result_extra0_reg[5] .power_up = "low";

dffeas \result_extra0_reg[4] (
	.clk(clock),
	.d(\result_wire[4] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[4]~q ),
	.prn(vcc));
defparam \result_extra0_reg[4] .is_wysiwyg = "true";
defparam \result_extra0_reg[4] .power_up = "low";

dffeas \result_extra0_reg[3] (
	.clk(clock),
	.d(\result_wire[3] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[3]~q ),
	.prn(vcc));
defparam \result_extra0_reg[3] .is_wysiwyg = "true";
defparam \result_extra0_reg[3] .power_up = "low";

dffeas \result_extra0_reg[2] (
	.clk(clock),
	.d(\result_wire[2] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[2]~q ),
	.prn(vcc));
defparam \result_extra0_reg[2] .is_wysiwyg = "true";
defparam \result_extra0_reg[2] .power_up = "low";

dffeas \result_extra0_reg[1] (
	.clk(clock),
	.d(\result_wire[1] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[1]~q ),
	.prn(vcc));
defparam \result_extra0_reg[1] .is_wysiwyg = "true";
defparam \result_extra0_reg[1] .power_up = "low";

dffeas \result_extra0_reg[0] (
	.clk(clock),
	.d(\result_wire[0] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\result_extra0_reg[0]~q ),
	.prn(vcc));
defparam \result_extra0_reg[0] .is_wysiwyg = "true";
defparam \result_extra0_reg[0] .power_up = "low";

endmodule
