// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
YQykVqWwqBHFheMgTC4RZ4CSmWun1pIcdb2fIiGBTtx4Fo8O659kKYEt7XfLaWx5GjIXFWYJ0Faq
3lUDZxsn+0AQc6EJkijszp5pbSfqIuGzP0jnxuS4WYeXHpd1byZj23g8otdm3DoThKqNTAN7W3gl
rMC9wTwiMg9UMRAXy1JOCffqI7mB03axXdTKfELBFv/aBKOtudFoQLI7lSqJTMiieS8bfsBz/ktc
QSYhue+B47wtnLY0xVWGKy6ZoKU+mbfWkvLKGT/uwzhZ+CLK4PZqHf9gytBHETLtGl8xAOH9ahF5
8sJP2LSTnx6bBoZnuYb8KBt5ENSARwWy/cknKA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 1680)
1OVDwvp2CANv/QoQuaMqqdnAMKv7LUdTQfoyEB/+fSXPNekancWJeCXycThu0LduljMbE4PjVfbK
+q47KTuXSPqYov7NHbLBd1EHtX0oYUi2opTLw1O2aI1zNlCXLy3GekUXC5tQpS+u+fkR6WADsQkQ
ko1gUkiDwCtyD9Lg/aMDEX6HEQMtVFIElX0PuJ7rIZ4ykEAdM/KqedMtfoqafn41gGCVKLvRqAX5
9jv3Rgqnk6maSjvzoKNRTLzEVK0tNcL8iN3ORSyCldkLXbVYB09WcGfdWvTMgLYbH3ry1myTZ8xa
72oi8SOTzc209GUlK3/V2jplc/74uCFS0aWVTjS+RWWWSKwFlSIpPgAmIrM5lCVud5vQnPEoedQN
U87lfrSqYlChUGYu2+3DXh4S6oQK9HQ7NvmQCBhMaZHeBLOmxOts0itGrw1a6e3M+iH9/HvAMArf
kcoCP4qVBfmnoVztBrDbzUBtIAitRt3p7b0GdTxcDpqa2kRBnsHddu1m9YtYGpsRQk/vQ+be2DnA
g+mRu/w25hrCB/xh6dwnLTy6kXNqY0y2KYD8sypw9q+AwBXTZVNGoHYQ/1q0KUcvHexF83L267bI
t1bvEGOfHSaPHpsTCHMVKjkOWqcbK7KLLprmbPMGnN5LC04HaN1cJlOuaIXA48k7BcPu3J592T2M
FTnESs/VzvgTL4haGWwVqvBpwRWkadds/wcTTVHF5d46I6MB0iXkFnyvG3zkfvPI39CJJ007dRLP
WkaKKKjgfK9IgDHkUsfidNuBL4yeolRugbColNlLy1T7aa2o+k4m4hp43+Ja1vYjx2FjCTcuhIxD
XPM/V21zEgYwnPOlzKUYu2+xcbex0bnxV2dCqjERjtJcJkunmNCcMAvJdjmC6xJtI0jvVkUwUg9U
2nO5wxZCFezCoGJ49pjuGOr2nyFz1T8GScF45YYEkNvxqJlShKNIFcMXcM5g+J16vaWAVCLMvuXN
z6fya2Imod+vGC1HrVJauBFwhKG5FrFCoPi+YCaQPMFpiyqFCY+SS9F0YcBJJy3icc2pCYnVywba
KY6kNko7hawGF5SRHJb/ZPJAGeghS72mfgQ+Om56+mL4vcMrdEu4D8CApEPYpUCgr70AlNL2sgO6
70yAUV86v5vC8uLoznxIbewy1yJwtbLybYmWLKHllFLOxo2VcxiodA9LkcEu9R/i6kuIFv/IQhVv
5IY6txBA+L1VI5dAoHszp5cJ+g7u1Urr3AygbuTy2XCBznj+Ch3/c9tdSi5c51VsdVihFRkB3Jbp
Vi+ySXqYlTKXetoDpHeKpmbiaNatFy9QUJS9iTGKDuDuBcupBy/FAwnbKxmjHbB6RM74ACu/Knou
SzSQBH3RUIxnRsWuVy131ckgH7JiDDanWAHPtkQtyqiQq9PAGj3T82IVv/U50cTNIzbxp78PCpBC
Lk2h7cDiTMOhVxO0atDkXAfW7UZzuYFGxCAUP4CCUXrlgioJXRZSsx1sDMJgtdhGUHUc8yrPx+iz
0gyHBztATAYae9t7MIHEY/22+Q6P/nygaTaJ/+0GuwLFV8qnSUZ2d3J7NxD94OV4Vh7g39fbQ0xA
7H9vkqrMzJGh54+VxflxxjiTqSdu0HCmA7k6T/1NPM0DKStb3rsZEGyNyd2O70Nx0kbtK4I4kLYC
D3VcDYmyG9cioEYxe67PgF16paEA2WxZPgjMImQICqmH9DOALFMgll3L+GXyXya5THylT22bZulm
WS4oX9Qg5/ypp+dNGlmF5r2/1U5bQPQ+IFWLDhRnb3IZXkhy2qA9s3KsOYoW7LvO6DTiMha23hG7
R9KuQsxgNwY2UbSWBLPgbQifwPEoMozopAB7cVDKuXPNmithYk7PO0Ytg+u30eaHrvKI84fMq/LN
ESaCF5K5cZSssroAdpkYSvKyo10oNy6mmIW/E2VW4TnI9bYkTqKsHehtrncUc5Rx7IlN6iI7ZcwH
3sWkIoZk/Gv/SWHxPCOZk5kd1v2GVZ7mFSsDnC/s/tqWX/iAH/Ac/3WWDv1kICFY3Z/FipCykNra
T0dRMFjKoJ9JYYljSx87OWo6aKUlRIGT/lynhzajwCU/APFRz+4aWQDDbc19sWCfai0BUoeXEVEk
NrtAe2xq39q9uoZaMe53Pec7dai/RRG3DxQ5eOKQXdVU7b6/83vlSOl7/pI6FIVMPw1GtOhVYrZZ
QC65FPlwTn9ZkN1dbZaSMEfu32vUyvAiKloi
`pragma protect end_protected
