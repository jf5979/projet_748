// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ttJm0LQTAnT8JgJvqYIW2mKUnhqyGWfqXKXgCTVRisjb5NFuAs2+qsjqGkxwKu+78t5pENAf8IEI
d66BJJsJP3W8yA2Rt/lnrThLCjRnEjwGi1jJaE8cYzZYJIb+g2IwFR63xrtuMjpbk/5fBPf3J3aS
CxmthHWuwVhkTdJ5HWsWzqEDOCI9Z0DJ23MS+7fRu8Nf3HYafGO8ZsF346IzWI0GtUo93LpNWYOn
BAynVLjiPE+f2o6W+4rqYXF0R9Wqw6bRmGSVgBfMYo4MrDvbRjApHDCJrxnoAqsWlyiEwTlPEVie
/+W1hgApWm84XP7L3doe/jSazzLJA61qX8mhHQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 30032)
yyoy+AB4x90UaLFQyjBsYv+9Y1C7Ux0KP5iEFRa9uoQwVDDkkE8Z8NM+FcR68xOnF7vZNgUvL3Kq
Ow8RwRbIL059TkKAG495u5UmDRSRajIxwWK8Gcyk86oXDza5e1rNo1BLnolvMvKKx2poFBnjGBe2
jRga2L/gFro1QVlC8VjZ2Fcv2X8jy2JLJSSwW3JnBAKYlDv8h5+1hahEePDdPkQGR9RKv2ywKi3U
Z/t6TPxxQ67Me+YmSVV24D9DbXQgMPDItKd+1Wp2TcYm/XAekY9YEDpTVOvX4pfUWOFXPby1BflT
AaHY0+A7sQI1eCCQUEBIO6+L0tBMs1ajHlbzz6Rp+I9HXElO+Eh5rc442XGV9v/JPfcAQEH13nQd
7m20Ov2Z4koYuyNi+5R9dENtY55CkuXlTnw+nzjiEypL1QLFDlArb85LyNfhHCXe62jqd43l6T3/
P7dB7tmAQ2AXEjHfZiTRjV9+0d07xWT+UdGFEWgX1VDJBxoFnrBkygleliJDxsPZy0v388M5jaQq
dTju/qRpFFqNnVX9MAUNwsTRsGvV3yddHTzq22sSpAXo7fqwKdu6ERdRVZwA0QIsgh+1GsZga3mm
MBxIF+eVX5WcFlokpsr4wGOXURrAJdwP6/No79q506sCIedf4QRMRUoMVo4lVs+L3vTn/85CjN7o
oEveujor77BNiD5EWah6Km3qa6LyUlmWaGdT5nzgU37oLR7z5YTKps80dLG5uPj5xUFqPLNljZTc
4u/83+oKRzpZil8eMUQwijbrI6Cx28qcjWQCOQXCPxB+Rkwel7KzBpE4vWfiZSGtMY6o6YAWxvsw
32yk/zu9D1eGNtIw2NqyG6fKL46b03ru/YcRlwAuKip+3s7tiQYIeDRG99P/3Ct0koj9tliy9bnb
lPQtFz1Q+ha0x+J02gZUMbG5wRBRGHPdtdzmSFvC02YNb2xdxFOb205yuh4dH4Szkfvt0YOYH554
sHULBAYg68VhLl/i5gZ6nQ+dRZ4fQ+YRLEcYhY/964aMqDWUqROclMzWAP2cJ5vlj3y24twbGda3
tpi1AazFr/INzfSoG/71jfNYy2U3lZpEyfbno7XRfzRKnY6KSfKKRvezOK4FSvQPmwD1f5bbO4Ea
mFNCcg91xR9cZ1LVy5T2XklAPx/gCX32mnlZ4NPZfp/IYtBGud7ZEt1hojpJb4MZYMrZ7ywJj4wo
6++d1/nLJgvy+Jx2viQ7QNjczD1zk38inGiSs3iQI5AVhBhsc43ezjIXGvaU+TP9CfSeRKlHENDd
WPY11Qgjj3Nja79AuGj7PF46AH8nrZqXBRbYppV7yfJpLU8xftZ8zUTA+pbQgHzgfJpCQH7Iym7B
1F6U8O/1SsyvEgvpfisYj/8jP6LbmkRdXQBHqAWrGBOtRq/pZxqsUDPlfgdDYAJLeDS3RbdeJvKh
ecOJB1SIBeW15JW5N0IFKkLBECrytZ09dXL7mIiqhFsLyf5tpxPdcpYRXu8VcKNf2doWTeLHr5+K
EDLrgh1H+BIRzvdGVEWharGhYz7AwUmNo3JohlTedmLrB3s7e8M+r3tFLk4FrNZXf8HC5DR22evl
VI6zm1jDdkYJxjUptfhK5Rp5d5qj84yPpAi5SpmMSSBHYWvRJ4ekCmzvxnGZUKs1KGkUCHtd2TB0
hvl2nJ0ymUHWWNEWk0OQ32qOrcpYylUyJ5N7zN8rmFhhyj76+naqplfWeDs/2lWrhJZEv8veUo/x
VM2Mdzk2wa1CDy/gKqV00xKOgN/EB6CTrA2W1SqOXlKS8Bhex1D3nCfu5vXVHvJkIOj0RBwJ5fin
k4R2OnliII/Oo8zsNVfzUcV/4fMsyhpOI7ev60TRVZGNcPQCAwueFQZ5it5BypYMVGxDL2BVorJb
EA3D6sq/CGe9x9/4xGTA5+qG/W9hwqzsVTlGNgk3CJMjN9D5/ijMhVEkTUHU/EClFC6Mt8j4pZ/x
WYC9+felBplOO4KrKNbJMqymUmMsA7X+hje7RxKlrShF70YgNOqFeB61PgjtjYyBgELZ374i5ZtQ
MtebSekA70hmDQZq8ihOzfRse4J/ZNMmP2F2VSbAg1D/zqMDIvcKnJVxOqxHgQ5jTtB/zxi8HAcV
WZsQjsIBMoTCnZU7P3oj/bO1SxFnjQLrz/xgagJljk7u7tvSXEI/NkDLTumkZ1rY6rleDxw74ibn
6D7r7tK6UVBMdJeXEn5knQYAC+3jtxEQbRQxnSiakaotVgoX+X0J3ORsf+5zfz1TchZ7t+avP4ZG
HvXKWyD1ToiFzfs7NAylU99Od6ouoWkZvdIc3NTNp5Kfkp5MjKlK74oU0sYlS8aWiMpbrNlOI7gI
iQf8kSVv+F03HGt4FuYyEh2j0O0M2FRQOZ3krz7oFf5fXMSEUz4GZ4NunVkL2d0SL60jOApbkQmt
QqfebRMBJwz77kBbruHGAL+Dt3Qlc6m9r0NbUdoWNT5YIl/PErDixomg7fmDcDdPgdos7qAK8OAP
6Mb0fur5hmdJ+3Agx4bYo/DNnw/vD6s4zMnltBdYoeXVnEQRqIBSLZYI7dieW2Vtj3jHY5h+SEEJ
NvqnqnNarJiwrgGcjy7GC+ABYRiERgIlC3qpEIqeBL5eAKRvRFDK7LNgCZ+ROvAbTM8ish2x67JX
59qOWtLuXHF0ARdNVkKOTXrmKqDGaWdwX8+t9d1FeWHm0H3kw+/LMNnBWlR/Nw++lSW1RV6djDvf
ueH6ZdjjimdXpBUasZKG3UktZPCgjYf0Yed/Y13iIvzPWIFuhaeGFuflK7jBXHIDs+nmho816N9f
7177t077hDmZJgRl8IIGnC9onZUTapDi5CsmDlgemGqjeoLFAc3WCRDiQp4JEMC6aAREIVBJsYCq
MEsMVHyFrxKnN++XWDHWuzxMv2dDaK8xDiqjAKoWis8ep8YHLrzozrqHU4VYYhbLrFeJz+cKnWGz
R6seswmaFoJ3NYfHE0jKJgGvLdZsO1Zi4ha/RD/mIuFAIS/XdvR1cg8xsOBHrNbGD2qaUcpyAWoH
L7HvQ824UcWEEPG215IFyD1b/knia3Lti1mOgumIpLxAGvbxgWUW8VMdEq64FCDhtHx6NYCa+qk/
nGs6wdLbaHP9/cJi4uzg2LIQfIWbfCWJF7cUvZ3JVOLeyeTjoWQN0eSwyk28Kj65/KP7l+OcQ4J8
0DEQhvemvY8T0iYsn2gfvPAe/0LrE7OFE7Fg6qH8YFJoGmgazxgIQGdjMWrBF2S1CwWcVrCUG8O4
zBbfZYeRkaGz1q0gmVJkkJPGqYkd2Y7yLSnuW03y43KpjJvBJgDUZkbsDo4n6z3H6tl2VnqasdSj
kO26rHNAuwC6a92eYM8icfmu4MQnKmrnBgvUI3/bMNX7VZrUorwuzj17ekLKFW2Js83XkZQeXPIM
4vhr7q4J/7IirEbdwtSJutiClJCyaLeb6lp2uHydMZmRmG3hZe+YHZIVRqWWQulUUPx/6nsd4M/h
KI/Z5YtiC+xaz63Q2BElAiHGMqR3+I/y0hOKMSIymIMShMilbWCkP0YMX08oSpcL6d/OW0LGAX+3
s1VlUL2aVaolCv4jNTRVHsF8slF5/PLk7G59frXLSsJj1QbNKNmY+0QZwBosTn8/WTkAhp5guyi3
porONiWZp5MpnPOynYuOTN4UWzUFoWLy7jSIDtTrZozn+yZ9oyhG7rWNiLdOVyzve6szie4nDnfb
klI9Lf4oaynzICrSwfc9igTDYfp/ZqAvuZwxRMMUxLJr0h+0tr4GJTxc7Bu3A8P7OzrlBllkDceO
FyraR1TXRt5+OeLonMhreYvSd4HYB9b5nIna1OUq4Rl2k3ui7/L22iEeP9D6BNLLjov4ADr0cQWB
alhMu4d/Max6XZ1/FQEq0TNJHKa3GJSSnrKfJDO/7jboQ3PLI1VDpnJaQj1kyf5/rJd11D9qMO16
5eEVEv/wyRt2De11vfYtzlg1h6gj8TiNASwgdCecXYSPabWn/MSffVSzFuSej47eNaklAwpc/6/I
pTVbMSvGy5vK0i5ecg/baBPVqrlOueW2PlRP+sJu5iG4JC294g+7nY3oVm5Fo8BGLITLzcrXf9jg
o+//2C1/WhW9sBfPx5OihsmaCxpn1cKAZoVInn/wpufyHiG12f4tT8rwCXkqLNhG2q9t0F7e4aYb
sb+BM9A2ynUK2c0/W44DuR0meBzNPFbwJf6VM+WDhx/VzSdWmOJeBrHqZZ5c0qhotYX8rhzCxHor
X1oaPFRlsm3OTY8DOfJY7Wsd1OZtiUhrflQJkBtO2oOJAReTjj3lhzdH3O3kgkQsNw8IS0xJlHYJ
p2bptiF7wQJli1VoKZUeo/Y8AJQv74uPiRCMZrqfdhbUL/1a7pe70cc/gXc724OWLHmRE+uxMkY5
/cZnG4JvBOdgEYMoRxfSmatKE7vth3YE4KNQ7R9AFZIgholRjVNX5zivN615EU7PGi/njaMpKqUZ
4JCcYUuUZO0PZd+qCU+VrmnONV2weSdatSTxDWL7uMxoYV1U/8zVz4xzwskysiEylGkYwsugTx/Y
teB8oaoySi7kbxVaQu+v4z7+JgnNRDmDud/v/f2cQUVjghKCgVq3UV99cMndJTJwumo9OOaljcRf
oskYga4yeT95+YgkWbX5kDWyMBLGobUXhKnNGnB22mC8nF06bff6kofczyP6FnH9YQ2Gx8/gAFiU
Y5ZhHJ4tjSmz/3Uo1oTumzrqH4yadRL0EM6IBEaKc2+zMWQGM38aUKnxp98FdSGbBSgS/YlFyQk0
Y9aLGHGv5BcMAobQk+UvcHY8KslBI8uKFM6y+8oDUz9Ka8D8eoqYHYz+QrSLOs0H2dAsrZVTw1Yo
dqNeOfTj+nfuhQ5bPjHrCL2JeGNJKZgvRp53sv86MY+hZ/bY9H4GprABlB+Gu06uWm7nZNRVlSMc
dXLp+qoBDiZwmkmGbRTvL5mbWx0VDqpue6yl2TysaaHfy+Lr2TR3BrHlZ7doOF/D4S6V1cCHCPJS
h1cd19MQxuhx08iQ7xE/UkZ511mqz7GCWgyLduL7/3MLZR+ZPRNeXYedde+FIhgeQiujIvK0vxOC
1MqyuCV/eKghZmx8oE2vdw6LrjDa9KCTxzmzHd5/IC3g0QpxkY0uYAaRt+cweJKs8PaWJmjjMLF7
1JCaQjxyRh35t8h1H/ZuMEgh0Bs99jHaDzDYFsF7FALG1+CUCH0oPDhZPK8uhtHc/+TPs/DNTIxJ
b5hJgONKQ8h73kVzqISxNjW+Rw+d66mvCtE0xQ07SGLwL8xedf6ZijOJ02U8qdxzKz+tPjwWUrNW
AlWMyqVMOYPVBxfHU3tWuBZUzy95k/+rIHALZGTWleDkcV68ob4YBSCUYEGP6DIRoFPlaOUz+cb7
pBZmz8U8dalovIaGrFVzD+JRCZzdmshiO4ye/NLJPBItCl+p3UJ24L91OVUqAtzXFLnAWCGMZsZ3
VuvSggIQZvNFokCjMGNJ4gvufCceiCbB9Hr097QLlOj1Cpdl33K/7D+f7NBhWfj65zsVJagKkI2Z
unqxKctknB1mW941m2i5I++gxjCsg5GY2T/hvZofvwTzp02gtpiqxOUN+SPoo3BLw5hsRRu3eksB
Byqu7cpwKJpojBMmlRA9eOg8SD5b/C4WbZtzzDJJuWB/4uOUPlM+O/CHgO7vy7G1RvuS0aFSmmTa
YdBvyZrW2SaPc4nAiueIC9pkJgztN9zfqP5Y456+xbQOaxKxUBPhKOYt59mjAE9Vob94CbhnOZJX
BZk9D4ZoY6wVgvGMB9UjeIzyKSvA44yA5g7TBHwSx707tli2Rwvp578wUbKBfa400o7R/IHcLOMh
WCNRDursIf1fXMY/DMIEjrc8p8nUz3SfprsFzZtmzuOlEBdLM8GquXsSXAeNrbqjLTUnDQHgz26j
6mIk8sKDVlhXBwfVNQvfr/I137KJORmT/r64t3CdbRo2uhMCbt2s7TlneijB6DQkEfRRgu5rjnj9
mX6GwypGmw52LQTuCnME6R1ihK5MxsgJDYKvZAuVcAFnX6uV/Pr+Z/DoGbyaMySMpvQ5pyCvL2Wq
6vtW3XzHPR7zjUht4s1He42y/SYxrcFSonrTb15H1nP33DOTeHNu0Awwp8nN6yLAMMQzu4Ohr0bO
U1m0UKNAVeOIvJzYaEmInB8MtFF7+R8L3rJ90dfvBgsXjStghFNslgj4SY90Hnzx6lK20SIi/Jsc
S+SJ/6FwSdwYJw/BU8aPNH3gtCODDwu+pc7N0R41ha0KzA5+JDxolW+9o3xBVJoQUnBAxsbKiFD5
kURUazsM9OLyXNSRCcsEJYAvjREPk6OKKxRgY5AhSQ8T6q6E3gq177Qr7BMym8Ri8gC1nmsov1AG
BTe6307dKdbZHxgSQAwEE21P0L2Utm3X8t6ERQhDkusUopRqAW6etVn22b7YCd2qH+S5xE/KN0hj
Dd2iRSZaIUwuamp2cNYQgSV7UzceUQzgI0SdrwvM7p4geTHw5SV4LhWKT5PGcKzm6DksP3pXNnMp
YIY5KZW7eyKCvOUfEl0kDrUPMsNTsJD/bO2qpWOCiIG8bQJCH0R6/q8FHUCG0GTVbrjbp8ezMy29
drki9U261cdNCllhpLbBRe6dISQYROHK9KpgK+b5L6JAgH6iDhj3uErgB2SBm3B2mO4icsSnwzh1
fuSFAD44Pb/31BGeWcZSjCjITf7y8b3DW879bcgrQC1oxAmgbCVyUqXMdWWyj4d/VVw5iV7x0CIC
6/+xS7dwoyRlw+wAvFf4nCFpKQKVR/U+P+tGEb3x0TISN3L8Q7fDP0cfZ/zNXm4u/Znkn/2L9GMH
48SmFr1XRhvMZMRjszyEf9mCTh4O+MFnL2i/dUMZIt9JerZiKAGVS/xdunD8+gNA7N+aVHayk/Lk
5MJFzTXmaSOWq+/Yvj1V1NHkxv1A9BRbWNzuy/LdYfyAM50nDpjX9EVNWAgERaCR/rEdyv9zSupB
N2Q1fjV44mDltQR2I0XmJRdMuy0LyQFdoUeSnUDwoLsl5hANG3I/IEJ447lduvfY/W7nOx2ksvbA
D4aSM3bY6JYIExWrMaaz89WaC8wL4MMiwgB6hI5Q6oX32ejKti0GjDc/2Umo36VywDGKra6Hr1MI
vqxIkz9AM6R746XGZg0apxH9GdI6EhiZTxFpDKRYQcxdtdWWpI4LAZscfEpCsisBRplDHgLx70Nw
MqkUtuuVj+1+126WeYA2EjOTo5YL8mB38fLilo1C0jdMhTmNGVKJxPPyFPT6c5wTT605cZ5e5bDi
hFB84/pFZT6IXdoTdw5uoKxDfm77G+XesEr/HbntoAfoipSYT1rCb3auchgeMTD/Dh/iofuU8TYu
Z9iOpaV4FYEPqAOHDnV1pBw0dIXJA1qXFRBmWzknQDw8kL0jmB/eVWmNeStXwHk+NSDsJEZPLZaq
fv0923quKM1djB7izqec4QCjtfz2gqFrAxOJCFOedMOxP1MUnn85vRb9bKBjwmTfkgCD96PRddxe
ZqR/K0/s/qSHnJCTdXwK8eEeDx/VoRWA7D2XArR8wXuPzQT/lN8KYmtTJTsc2yGFjmkW7zjeAF5E
UoyNGmH9lu5p9TTZJXivDfSu3Z6/CQrSYv8WwpK6UdA3HuW5P4yRT5v2ho99AkndGlENkiXWqr6J
krfoZW05E5h/IuTOfRxIoLXFwI47EfQKUoHbNxwbqjw0ES73LAsl46SAeC14u5uZ+Q4Reqk5IJjf
WH9OxMcU1hldq5y+tUF070fyPTP0RSTeBom77W/FYFkOy24cOaWsAcrH35FeAqf58QYOAlnzKh36
70wFHrcWZTTHdyKdsl1xWBhcKUmjNNARzh5ThVAjw5IW+1y75UD4NpoDWTsNTdJmm1tN49tLP2sd
sCCVotQQ2khUZ9QVfVhvBowUuJRP/45WMzzftTlyjum4DVIiQOWbMMJJNsuCrangsDXRqdME33R3
eq/t0J/XCXnLL928a87he0IktOtvtI93IRVk3NzQPbEmI+iv5LJzp0eyPKbl6/53HgYxihgxqihz
EtDxpGbLv0QkQDT0iLbt7hoKeAY4kcjxhVpy7JjRqLgSmECTQBq1B+3EnRQjJ1/guN6+JhXL3F7y
7iYNUAnJZFI8vmaQQkA7LIfJOxPP+BZ2hHuO7TgWHZlavbZUugh4ag70vnmEtaSHcE6E+lPda7fg
qMJ85TtBx2RbmYGw+45zA/nByksANP7IqHOsGJRoEPb37ws5sSrmlOjefwrwu1sn4qoTQ50iQz6m
x6B7pL78ftc8pa7LeDMcNs2tnR31/4cijDrCn63/WOHXNzRnvHitkq8XaQqhqIqfHHbA1LNQ127p
N2jhALpFQTU885DNMZaINtdygoT6CezwDLv6nxqo4JnIzPM5BQ4k8s1Qo0y5uH2bCjBXvvaUNBWS
UjxjXwJ+BLv1NluUsnaQc1ZO6p8mcCBK5M/LsDDEfO86yjeePAdMVE8OVghEP/KD8CJptNWhOuFq
GuKo8Sxfbajm+ByHVzEDw/x7J5igue7XvmomSgXGWG8Jw9IAYFXTaHvq26tHRCSWxQlOgm1v5kuq
jqGgf6LqLqMt0vN7ygc3WUfyFSRQW/ii0auLrzlNAzbLxlY12dXXx3OYdkNaNTfFWIMVa7hNG5MV
nl+TZl/lLjxtKvJl+O0RglFpN7jYGJb8kk4LvZvBa7BpJ7GnDJ22FboGPDoUDqThIqHZe05SWHON
j6blY3qb1cYxjgvdOmJDn6iYI4tL/0PYc6+hHwccO5cHOduzkCufd5TCpIvmPmYVfST48IqkEilm
2Bo9AquVwM+8tmrFicSi18Xx4tStts1GwFI9/CWyWWkTrnEAZajoQ+woe+/mvMzpMNcQGni5IOyq
hi04P7YAciffBBBDm0DEU9A7U3LGyPLth7HA5cWrtBn+PWmqWUesr3r3Nsg5fSVs/WHHtmrbVxZj
vA17KIdHqJvFoFRGEMlbpwC2F7wzFH+Ivmvwh1Bf6mRodE0Avap35PLc9lRiMeuoQDpCxO4yztsd
izOQb517+Wr3zOlztrevMEyTl9D8HKTt6hMU9k8L09gKOpd5Xvf2hAFWhGtgAcovbjDevlmpzWsK
cKB61QyqIDANVDWzXqn8/wj/tYHsddMh4QSWySVzcwUgrzo4LJqRYJhhhsDQUJeWEWkkilhInI9y
LbO37n+HNAOwftWc13QiYM5jxK9+gnxVoDbnJgBYdcEXI1Vb5COsY4KzXvleyngZyWXvwdwRmBuC
uDe8nPxuCUVDVqgBsuT2+TtTL362icEqS03ENniMiF1Uur0a+h3C5XXz2B2VXM9w865nBgasW23Z
M7dTiIHmfj5CaqIbRhoreFRn+WK8NiCRXptngNqnI6KVcMeM6D0ESBsC7CZoyac3SOWWLX2zYUl2
cWM0lKTmIJMIC/gUupdQ7DrI0GR8SxzzwgvDAg4JeA47k1/q1sxVaoz0MQ13+MTH6PkQR5I+vHSx
AcPGrXU76mqe6xTWvE9u4eiAjJgwIBncaRx4acdbIvxdGNJ2PVuc7sHcoAQtcuwGjIE//xwdHU/B
aK+YzMh4SavoyfFQDBwYJy5lWXIowuy/shY77xT0hpeG+WxQoX1XxBvFE53f9tW0TFctFJOBnd1Z
N4JREZTCowFnqinAVzcT30y1lqnOlW/uIhri6kO/XESE/2xaHsPmQdKY42xpGwLJ8rHGNn+1YBl2
tZqK5vE3qk+17QxHjaNk9RGOx4snQVxqL4LBrvvV9YEepRr1ahdKarbtCgjGH46My7+M0vqCGIEP
nm5GtPyvOKD1bMSRMY+ANUqQHcbhuOEh+fTulUPgO8d5ROPk9xb3vyq8q20OJf6YqDbfwmNFOANt
7/S9lleq43tpPQKKPYQfOA0+SxCbZJ895yxkjo0AqBDuIUwIFGBej37mcPaXdU6ikRu6S2kDcfZ4
kysO8MqWOtsCkAt53RowOlzmhiaQTBHtH709uxrmMWf57vuhAseUzhAsnc0hwf5CYWJl0gfh6Qcg
QDxbZQ2ao/O4dD7w8TCEzOjeBcVK0yo0fw2xZg/gzoV1pG+UmZl/5n+D6BFAL2QbzfPTrHp8ZXnw
dfs6cd6BDGycadzAzljjtJldEtS+s35c8fgwNKUrVfjzjP6MMFF7i71xISaHwhlqky+VYqNUa9zR
znMhG1pMqRLn9qdK8fnxcp+ZBCunyX0T84KtyqTyq6BCpyZw5JoAQTGyGQTltpv+Aeue3rewUtqk
4xAQO76WQ1jlcuJh4Fn4oXbss37v5DkroLKmjDfCZItbFeS60mYnJUxmfmDlZ8XTPNvf5sZgxsdW
FLZn9+LHSeMPuzDPXazrEZAfICgP4Vmoptx4g6IHlA1AIht5LPuJPKFUzHhrt4gRTaYifYvC7Q0B
0C0tBW8Ke2Spn6vaww1qNtXUCYoH6TFAtbUtpN8A8/LxtLUdL0WuAMJaiAa25m+NDFQshksclFsk
ieoLKZQCwyUDHw2sIwuKHsivJ6ud926tABAPlbfxV4jA14PgK7csWLIbmzAFMsf2bKtv8n6o07uR
pmgnnwfnOCf5Nw7JSmmLq4aeliQiddOvtdOpJO8cKjw65gttWGkc5orZ/94eXrwnvEtBZm8gIw0b
avtRK+MPiDuqHgjJHpOKm8XPwojFrHSmHpkTHEs6dnoH2VYKGQG0ZmvNVd9WeDr9raajQKRHrc6q
ywd5E9YqTzwmgKwRU23p40Hl2aZdwQph2ZlZ/AL/nYF8ltPBr/l9WoKAkr2IJvDYV1Ihafc8bauW
d4yaFSnn3L3Ns4+B5qSDqvO80y+U6KRy3EfsQRCtoKdU4OQ6DY8qruHhdYdvHHrRcA1T8hA/H5fu
6QFbdI7O7GsrB0NGWd1lef4q4HoeoY/vJHpZutKbUXKUSnRmJh/ZJF1qksvASMBaqdlkrcf2bwaV
xTIGoxcphL2ZipK6/HjlAHC0sDHpkXjF+cGLYokppJ6tzcXGrtMh/Drk9uPthd7wmjlALZyA2zm7
/sZlmttIsl6oJBZASpoSZQE88yox0RwoGTshEefbqkLy4b96/22WKXdcVulEf7l6G6eroqtAAaJ9
mPx0Aun2jyjsJheD54A4zT1hCM2OV804sDdDiULniQsetIUDG8Q8ntRIvLoIaOr9uha7dQYUpTw7
BfClJP2aD1cIgRbpm4on0WrYhzcqjpxkwkOhHn7bZ+hjVk2f128M4wHTSsE1bPRz2vOILxgiI1aE
2BpOtXgofXj26TlDhtvOHwAh0seH2oDcL5xqNGNHNv6aDi/NS0OFtPvbpZywOqSyjlf7JkDh4ZVo
PIgLeqpfdYJo/LY4Y5LexqHt4xarUAnHL3fobGxlHvt68Fi9L2QvTOAX/eDqAUiPRsPv7BF6k2aZ
vcBQawsygWscEdpkFY+dpWlHdL8gCX8JaccsBhyQuXH+yQejMYwiinMwOajLS63aNDa0KtW/kIxa
x+WOip2ZnNTIRxKJM8XmO3W7DEW40ZGZZHxtQSqgm6Zc7OFuFGU+NbYTX0bYDnWEinvOgM+jJMH0
desusI6E2wSNI6JI1h4Zmo5Sp0e5mfkLA4ZRxLBxPkm1JmCvNI+bbyiUxS/DP6LKFgEh4jPu985/
/0W85qfyWVGuOr0N5xIT/Y0qGkas4DvuApkYV7ivNfSWOf0sHZnR9ws394LDhFXBPAv3wmtBC2fy
7Mdm1QR43riPBMwTrVrVJ+OVue5YYiP0io+YGNy2j7n0ONhnJDwhTJ+IxPulE4PsWqb14RctQfNN
gRQsanMysFPADeX5DvhgrR7/9+YIBt51fGOD0aF1yeTFUIWmXWX5oh4IcrD3cQ5/gXRly1kDaI2h
T3+var2rb+O9iry6sU2gtJrq58U1haC3sA0Oa9sj2zYJ+nC47d/yGb9WzFkw/5dMv+VhXhfaIbE3
52AhBO9RZlFiso4oG/KKDO8iawxZ/EvtE3ukb4mGihN4N9Calp8yFEljWhnuDlagTaLcgqjgbbka
p3zL4sGu2H7C0NeE9zTzRUdrDHwtnfzUNYEGPe/9Aaqn5sInjxFei24sJJZHGTK4+vnZVuylJ2Os
1CjTI0zx0n5781pSLKpnqNMh9Rrc9blAUt/fBZnjk+qaGx8EUcPxCN+SuLiC/JAyhREMPCwm2e8A
fRIdx8I18xevtdW/sjD6GavlDhFItouXPVFhAfwfh7zQrBDDgnSJwNfoJ7r5rHIQcmeDt7q1b7oY
LVJROvuDQiB8YwEBMBHivyunPd9/ZCyVPqF8GG57TyaZ18htlh9sKsMnG2iO2NvhXtFGo7xZcDlK
FwAiuH4xiWLOSWHzY6cbtnHL4zDEZ0B1gpO+FVHZEQhbvO9JcQA+LObF45ZSmIFN+H9WK/DLN1YG
+euaj3krTvYQe7teHHlcTSlUc8/ELy26YJiMjDoXzitQnvivIQrjap8supvzAtmwUqPxMR1FM1Cg
y+2XH+5MOqPcrZviVpjZiM42Ikt1R323/Ze0Q6vbttH0McWULUaSYAKFMFG5T9g4ljmVlXopKKhF
lxmcACogBRIUaQV/Emu3+//Dg4qc6srtcMmX5HD60gtpAEQ54QCvAjEVw6guKC2R6e3rvayJEuYq
VaYYYpnSLBkMq5MCKxhsJoXuL7RZHi1mZNPm4xcJUpAvs4KyoAm2I8ZqVRs18TTWLbBY5zCYtcPM
nNFdxlAB21+SElCDBrZvLOG22zidDwAkpG5vOfTCqizOGJdE7VBJmndwiGW3OP0+1Y5suNYr1xvy
Pbau2lG5LY3loOeDmc2CzD6K9EK5ffdhoNI1kzSNguW6KLBKB05JNc9h2zxReKjmF5h97tL9utfS
SGKNQPcqIYdFu5JsWSeoMrI18N/+ZQ9X2OD0kDP1Wt1C7Y8Vqf+z9SRxi4/IbQAg3dklRi5KgjIM
y53cDLdSEHoTuvs+1Xv2pgEk1G3y7a874ZINxZu7iwugosUvZPbFRYJ9K1nGQkL2DEFhveVHIS30
mcp7b07qHz+bV5jylYvOaT/3tU8mcbyoc60oSUiSfj2/dqE/pwpJz/5RhTQh/d1dADFRwrpth8bf
u+Sldhb6IsbXVFjOYi04ZyW98NtHCRgWjvnE1hcPn8oLI3hixmMq3U7XWdtc+8fSNA0m/ztANQBG
QlFGW57X3kArQweZlta+uQu9oSUiw45U/PQ3eiqzBl2NCkCTX8/pZ1sOKYgZC451yCFf1XeLbkwA
vr9h3Fk9VCyej75QU71ktvKkaUoOnphi8PJnD1uc02S0+4IdV4u04SWPrV/tSthaYCiUHs9xE3/m
cRTBS5D93Q7u9xTSE4yoDq8mVdM0ZkWSVzgchBMCHI8mZz4huURotazDWZV8l/OJVouVufwPJDa3
3N9JlYMbK3SILGv3XcCC9Aju320KhDuRv9q9Y31cD1GX4R825fV/ZZ0MksqDLzF7EMuxZgLVRUmm
QsQdJ+X39fQkR4+c7PVkquSzzyG5n912OZieOXdHEEhuqXX1FUVCH5MQLR2M50t+KJbDyAcuS189
PlkUWyGOVR/Vm0kSQ0YW4+v2RSywh1+g8e1tqQRNkW1O8KQc5qC2+fU/i1P7rtnPTQp/47Rqr56i
lsc4e3oxT5C2OSEXkZR4XfDPmKgF8b7z+FQ1hG0g7Df2ZH7Jyq9Q9+5XLies+Ry52v+bjdMkrkVh
5sb9wnCT2K39+aL/AyenAca0UhfSWClo1OcK7cWyOT3p3b7faUCKNodB/lGeXNaLZxlLgGC0RQz+
13KaYMltO3Ofpbsh1W0ZXKO/FCKjwOkcCnYlHSAS07HC/7n92VGerxOI+AnjDjdozfb5J1cpHh+f
ZMKVDV9p6HXny0dzszCpkeaQPZm6KR/a5XMBXQUApRk6ZsNnQUrs/zDlEt8d0159fZcJciVJADMo
RfViJmOCD/SZiBU7ili0xMpidje9UKqmyTsp2bltG7EgE8Np/k7x/X+dHGJA0u6BweaCtAopVQga
ieAOPEIGt/wBh5lIkrLwAsDNAhdfSP3Uq/tsHPweRHp0Di34okgrXlRhqR2hfb5I4DfYlUBdw0Ns
DFHcT65scYH42KshaP6f+0l2Zy57BPr+2lzfqJQR6sLF/Mib75W/Vqrgt4R/88rBkg88Los6Qotr
eR7N+Ay8r5bqJZQmPHWnpP5xIfyCeN/QtkeDb+ni7J1/wpwCsEah4hkJXXf2vclUrNHs2YQmGuod
+loxN9ZP+QFuzq4UKD7tH60HM46ellL47RPg4qvUi3yDccpdUiwMaVYipLqF30sw/DKOBnc/Ush4
YIRW4E2Nq8fYgfoE9KdJgPcPhdx5rCe9ZMSFHdxnaDSDcJNIbYiD/ireNbDnF2HVEdy8mK+zEns3
yoik6JudFkQXnDO3/A/E7FFnxPd3kjX3l/sMZ+Q0Dh2vPWmu/osp+8GM/+VpwdDbIt/S+GYgknkq
6LwtZDr3jnEpWwtSnsfAs/8SDcbFj7kTvvBMPgl7AKei4Z4f9ld4dEgltleJTWMVGPOj5UfDZLco
+bHbMnAunD75eUfVe84rey3dfgH++IOwjcFlt14uyM0G0C4fXt3+T3ewUtIOw1UndKNtQMBURUgC
xxuSD1jGSf+HyjhpqNhA5OQ5z7Df0uKErEoYE6ZgMv15nh7u5TrJses07xk4o6uahsL5waMOZpYM
mIZVrwTd4ipqIOsJIi0pSavil701YBf9unwY5htEJTwJb+8j3f5UzVBxOFB6fW9sR3jrY1MSY+Sj
fdDmfmTZEBV+oydfrZ1f7FqHu1RYfvcwhAs9Ft5eqGCzCdnfU+G/vkYelgazygQ/eH0r3M1kNCkA
j6BlQIko/XfVDL1+umAPX3h5L5EXhQSjkBW6M5+apfgF2R44DKjqVDn1Fcevj9V6JMOq8ed1eHfa
YqA7OViHoNPJQkK67hQVsps+rk2TgdR4UerBvvqi4zxJ7qshgQmOxMFqQh9K2CcO18gSjYHS2Dre
CJUrefV3nfIooSvCwZ9aIW6+BhzLqLJT1Bs4reIQJvh3mZNm9Z0imLjeGvexRPgisPQpfwbQKTSX
EgdiMlitniXLY/yOlRJmoInBJ0yxA2UqTGHWP9/2YY80soMNwTH8RaqOPvHeTgrfm2xwjfvUS/bK
929s3F3yN3b+U++AiYPbkUO8E/27IFxrVxaE8qT8GOT+DIoiwS/3WD6dgEGkEChrsgxt+yYl52ND
yCATUhsb2YiYEJXjFL73b/n7qJnx92mcdR5lSzViS90/O3ntzpje7d7YnkIfTJdosxaW8sDS38cw
FRGMC8yPp+oKcLVpnTmDFC/kFgjpM9wbP9VjwbTkHO1dE3hxnHeD4Qodkdb5pwZXD/hKtR2AFgQK
RYuNk24atj1wERaxSLFAGwva1xuKb3gtBRp6aEj27EHm/twIVLchEfEr6p26WGzuuG7W7Ly5sSJd
6eLUWnTG+YeaGI0OP5SaC5ByMSINF9e0ISoduSJAXI8NRmmcfhDeiIdgy5Jiiuaem5qJRO2VMZAn
MOT9OjAInW5e0AbafLoAhEGEhR2V5iKlGUOUnbZWW31iZlxfGEu+qdAvrvn4jLluGPQeQIhJQnwK
qCwmN07Bn7kqXxqh2s0iNrqVe+OcV0cXYAv8jNCCqt+9dem8J4zDe5DQg43Saycuw4SA1n7d/cMb
oiI12IsiHghexYL+K0ro4EjxpxyvAd9jrlYWI5r6jN7oj12N7Rz/uO4+HsCW193v8zjK5ECFUlm7
/nwPciZ5IT4VL1/UNiRXDeCFMOaoaOrSxGkJlUC5ia5GK3H23jrpS2ZqXJDV56YcgGWJ8gkws7zS
WLSOsIIeE6+DV+y8cjG9l4Mj7m/wysnoGfYzR0XvIcywnGuCJEe/lDoKd3oY0VSA6CmH8dSDyt9d
/yZRUWq5INNW+9XErvU7JNWpNYP/QnV7k4aha8aochxD1DTmQZmke06bP+1nZ1CqmH3KZaOqqIsC
nT8BvPxDe5wXmLSdzL+oZLDVQ6jweogfsXXTuIBJ/ktDoqAhyokJWn3bWH76+DhrtUoRgKvI1fFc
jcNIfuV6M5kwl39kXKlVcT6TkjGdZii2nxxdQYqfwiBmkg9FTqmPHclpwv7cU9lo4NhHJ+h5HP43
hg7upmqmQJb7lu7MMtJ1oKdPuQgikBW+ckzDQeHicuOqk3QCD5XIy3N6gK19pUSI2JJG9/pPvV7a
ss7BOEjCRwGuMU1qUK+CaVOTRfYkRi7VH1gkn2ZpvJg26O+I6VGPjHtmp8HaUY61iu2lEzLGue8A
6Z8bLDTmrq35Md4p82KanNJ4xaNnxf5KzmgErOiGzqvGtiunJ+mAtqr2apTIx1GvwNqP9eA5sEYD
Pg47ymtVBgWxwGYiCQXl4X9ibdOoDXKvtb0XDsaQZCf8k+mOFkVTS3uaSFHwxrqlH3BCql5jgegj
IZ83Ionvq17mDjD6wtgRYv0K0GqXzoikCiohvBURZCY/6O8TAl+3kh118WcIB30ckzKhKvnI1xQD
kmtzvvSfGxFdxkI8aXvK10+k8pma9y0I8dEQkE2uiKqI6moTZhJwIX5qdaDVRZjuxNlCYguvN2xy
D1p7d/flWyfSgfHyuCDpXDv6gt8Ghl36tCTpjMbIzIpi5J3f7HDRjS/YweUTiI8Acr5AmJ5qGKER
TCLnff7/36ER/uf7lRe6nF3F2AwJsxPxozeMMDvbugTJMBXY4poe/k1lGW4xukgvzxdY6COfT8Rt
nym6rTN0MI0w4h2D4xIA7XoWzQSn+AmwDcu85iIQQeniecolcoIZJmedNPlBJNNGgnVZbgX/Jiu3
ttxugUqvuDchIbzkVf6WpQ50Uz+MldwICp0mXqTcrsH0KM7O+TRUendt2FL4uq7898jsbntcW3X6
Ckg+vBSv8hFovdbYdhYbYYSOT1pnyLiYe4mlbTNIKzsnpCZBFOWvvqaEdT6pzFUu0swN/C6N25t1
XFt2Lpl9y3RKv8tGgiAkPr8smlxCXOYwjn83pKPJRXpruZL3jC4HKpATnG6gyjqhxxuUF47TD4rA
+6oFx7CITwG33Qs4Gik2j0K8XhKNNqnIFPRFEE55/9R/7bfBB0sR8XZiV7ktqjIiHMZfexBTXq0v
rqpILGFBwrYNROt+TSbhRfeqYK8A/z5wTwz1GlrfG9jzC5YKU5O39HIBm2YkgbRNOe2dw97jLsgm
SJkG5yW0sXj1lAS+jCIUyhYFpSLxFyKNP4pEuPKFd8uSpVIHuddmtqO8mFrrixjr6fHDgGD6ZCOQ
hMqfZHvtcaONbnbB0+GGLCkn5Y+D+iuTaLmje4HpfDJ7nzmgcaWq8Hu2RkPRpKztk0nJD0s9NhYS
nKUAxZUEU/cLirHLdtBOtMdC1kEERQ9wEdPeTzDl7x6ES+zK1Lcwjnsc+NhyhSKBPUVzYQUmMbGd
3GkZz74v9axUdvYrN4bfkOxYvIT6+U6B23bjWkPHDM+RYuH99Ei2WbUjghw354Er48b9l5eZH0Xw
cZi6ecXkl6Wgdpx6Paqx3cPLn1FV2emZVkuDeePkIgCCypG9iU2PBp9Rm14li4kuLUnP9rSFnU6Z
NBYqYc8AYmH1fZ6OkDKI1hy2P7vnrkAHRAX7d/Tu1HBsl2pslrg2we+1+cn5Ontb6PhpXPzdYMrp
ZavaKt1rGHrfnsByqO1eMxf4dMd5JrQcwc7oimW14IIODkCpo/ujPIXOvdbPdVnqmz1ui/tZfKip
xbM+Ljqf95EWl+ziywkHWOcwtSgQbYDpgHPWqrCDihLw2xhwjPv0rxTgXtMm2vfYe/VW0zvNd9dx
2WFuAMg2nCvUIKSCfrbBCIQFSsBHaZ+zPYGP2CERUH2yk5nYsgizeGxzEMQFPIqcngjrFG0Q7hUW
KJDmeM0xswXKrDLKfNwVyiHKDVeXtX9jYX/YLxX4ptJUQLCXcDOJo9ymEnTDITeCYLqRthNzJ7ln
ZcKxiKmevA4PZLq16c8aO/RPOh2LlYnA0CTv1725E9xHjJzS7zJQQIJ37OIAehuHfJfHrLcERLV4
Pm7j3ijhx7RcjNqBWP4OoX22k9R0i27fQ3UJBpBVkEoxXMEF/I7TnHiGWP2XXwp9UexZPXJFU7oV
2VSeDe/LFGbfr1/fBI042gTbcEK9Yvb9RbfHVDjQizZ7nzM7WDEgYVar/G+fWAhMe25cQbtqd5O9
TBaHAnpXaGYbfQlNZaKBCzT+3eZJGzW92bhvD7fKiFolJdDgxEcJ7nvjn949unw/LLswEz0tsOFV
3PgyjdkTtaHTChsK7kebt1yUne1N5gvukh4i8zLgrZpZgzdzowaWRbrUlKDzUYOesVJ9kg0ks91+
49UHKxCkc1ybCt/PoY5syfYnhuZUWG5tfc96P4hgricsPkaBYKFz+uDabCFuv8nNSpe0laVQotsu
C6m83cqNq77AqkWdnzLpvJjZDWkpf8bMOhDPJjg11ZsckNuyE3xC6Ps4hFuQAflQBiSGeZlvV7h9
WArM+ZU+kPHz89P/FBh1o3sL0nnOVxVs+HIqnvQcNm+erU2/N8qkigSO2U8X1Am5iVA2PGnDzoxj
CnpgTjnAzSQmbxPi5SfH3YAGzhTZt827NdF07EzuzazLjshWKSfmXwYjAZVf4uo4MGhyXh5J2OwV
nG4BAUXgoOhDFNLiFEi0tXEHjIehItxhQv1b4Zjp6UxsUEiWGEK9jO3hO7OFaVv217NP0A33HMUd
bb8/lZH63UXCS0x8Cu52jtVoW2Tr4w8fk9Cw2vr2T5/TVba1+TcU/wC0pBqzibg481kKeYtGiiQ4
Ao1DNli+Q3D+8ldhttbglHsoujvqltIaMl4ZcoGdy3FKZ2fqJkyI7Ppc2GN2dIbpkoZ/pfEZQrKv
sU7K1XhCOLXuEPrVCZ4d3foqZZO+HbbAtaDpyFndOx5SA3ko1hyQj2wRvafiv1LZ7vRFXRgdG+9Z
Q24aFGDJNuVx7PRnG4bJQz/w2fupPHJ/eA9RRfBqKaJK2L/dC6kpR6JZNYYdD3AoDfswYlnmid1j
zBa0g4jrxWDDa5O2K2jaSrzgHarC4zVvv/mkwGr63QxaNR1/zrjUUARtYDmIULAbyhquroch5DEA
3d7ZJutqMzB6pt8a43W5MtT3NCXvCIkNlOKkhjirS1ekvxSIEvfQBdPB3e5bGvkbIjYRqePfEvkw
CEuoHgkUoIXqdS8cxYKoiuLV81/amdawu1UotJclrZqiD3VXLac/GaDLoyURi/Jv6pcJNQr2qFsQ
GuFE3VAe1A/dekMXLKfPNx5omxdwfLeS3SrB/1/WjjYlJ8Bw/UqQZyAbjz2dt1viDK8fK+J/31R1
j2b2zsK1Nb5MLCXZP3tEkdDuNHiRRudCdGpEHO4NqOy3wUPY47eXxiKTEr9JbXmCDO+WCL9kpNi1
K9PcpZr97XkEseIvyOmloibtbrLoXbLT+r2DSRsWVy8fGYmw2wooDczY8I2fphi6MHK9sEjU1pVv
C/atd8ulDHM44r+hm7YswyEjzMD30v0tt7Esssm0siW5GgkJTKzDn8zhH6Wg7ljeswMr0FYAQQ/8
LzL3vn1QXk31WhuROIQtoAiavcwFwMYT1nGDGURUTj0M4AT39m6X6icxyIb3ptdR5Bct6WfMZOEO
6hzcKL9Irjz8LSjpg51ix+n1dHQHSc30MiGZLxdKNiNsLzXjOwUCx/ifmipBruIhyYgxt5+CSI8u
FGtcLTIfUJdpmHXXXTxTIcL5ZDa/5EWPBp7eJWguYfW9zN61TgjzVzzI9OecFOcZPgEzpwhwDaOu
ZFYeXoOpWe3DZLkxbrJgB89/MGcftI9HViUGmsyFIlROvjwzpcLHy2lRsPyD9Ol8JaBoqrxkHUVb
i003Yi/5cI/wHgzpqvoE93TqBUbD+VIPPc/HE8FkuD8RsetEUZ1af92ahSQnXGxF+/tWkyTrmFIy
fcNj/B8sw3XFJ3ctrBEuwFayL3CRjyWEDVjWlMszIbqDCA0ou7NJLM0Y4DTAhIjMD4MXIyNYa8XB
WV/651PLtWqsxyVD02xCRcIqAgDsJJ32FVBhWXbmgNkExGQedDrIkjg9X8YzOMA1LaeglTvLUl6O
6C/Qc3cnLOfO5M76bawz8+aNdfmAPou0cfh1O7TY6Y1Dd1HeVrxCoRks5951/aQwDsAQr93W7JMh
80CnP0YE3g9pXz+HBkzIT6JnsawaaE1MElMi/OSzGFxIeBkSOEuV+OqyQxLsCetbGiieqz00Cv3L
F9x16h2a2SzYOZOeepzwkeaOORZc644SMDuTdQ2ujdsX4LZWY8/Mp4oMNjEBo8eMxSezA+3O2rjG
MTvyEFIVjvX0L9WYsJTRj0RRX8jq270KuDTS5niCw+Gaj9j+/z5F8nyIjKrh0Q+54gEJo2Fqq0Or
goC3x2jKHqnb8du58FrYY/Tan4icwDGzNPu99SHcbm1vND/e8QanI0JUn2xnuzT8Acudg6CCeMgS
oi//Z9hlEkFazZgRYgXr75P5BvBAXfXNTn/Jdfzg4ZN7JR0FRJSw8J60v59AW4weHUMwNo7USV2A
uaiiZilVvrj2bfb+SU7P5ggW8FE/1cOtM4ZK9x14soDQfzliMJPNYyNlAxBQACWX1qNssNYJa9cJ
yEl0BrPeqpNr6IiWZpM6XPUhZV0NzPnp++pyApwD3LOORINUbUvnkJ5hMOV/lGcGiR8WTOXSA65Q
YOKN/tt3TyzBxAaOfXcjsxhZKOwiv1wPytdu4dE8zZL1qwhA/E5UUkiN6SoJcRX/1lDxVVDaN0+C
ogu7nbeEadHQgK7ZsaxTVXaz/6Q4HhuzPDurWn56yy/Ioe9Bl5NoebWSA9HJ9tD3Ni07dGm7B6bF
N3ac9pGnmWDZsnmUKtSQkGhMu8Q8iLhUkUgWDNK01kHyPzk7MtXoVSq9ZmfPNi8pum2H+dFY1F3s
hMgO1x8uMgFNTezd9aST1DnvVKSJWUmBI45wprPqlDEDayz+D2H567E9SXQovVOc9upFDoBpD9Au
SWQ/0CQ8emq/ijRb1PjlLb6IbzP7Wl/37BhXFpi8VjqcCACEaqn9Pb+/bDzJn93ga99SaXqoUbrQ
0V/J1KOmzFFaKinQJzG695BIwWpMVGPhDE2G+2tfjVTKocS8WlkwfoJqyblElUwDDtz+qEEe8xym
H1SgMlidi0U27iVorzxmrLFjEMgKicrTj0wX4/8NuLOewjeCEVLIEOrdJPmg7RiG8K1HE85Wy6gY
1eFLnDFJnOeMndTWhWzc4HcRqYEc2PyJOvk1Y26oeECVcaO1yoQSw/xr7OBoYuK4a899aCQVxyJx
tEe4YgZX91glNC1egVSkCpIAnxLw5kJjJIW0/zZvVMyOlDoR8VPyqxRv7K57zdo5n8M/O7Ts6tgn
pi0A5LbietTLGOdZm+LjDYtlheNO1eYcaUpnxq6xg/mpIPbau42NpKAO+UjSsotzG33MP0V6Lr2H
PPYD21zJvNZLg7cTVoU0INIzrLtP41S6gs2JbdGf5ZyQmL+ZJ/x0mPruHVItAXoBuXhtNcWdC6/P
rDCQzg162q7zybKJWfh8rYDJfxaVZy+ATD77qlgqgLw87wQJFlQ+7O17Kxix04PkpFM9lj1fnYIF
mMwekhetjSLC1iUw8lORLZrLFIxNNI8ZSt4jHYldt7ebRHMi1jFEJ9lCM0vVfkREOW8EbfkhI30c
wjs2vngWMVX/eHgY5euQWzPAZdnsCr1qU5T9AN/dQY9/eDvV2Be9Rine23++F4AZ8GYhAbK5qYwj
3N1tB/XWvUYAuL+nJv9KNPKqkaEpRDN8ozz/tlA15ISoWUKSMwbhAn4TBSCtBYDZzpKAuz1vPTX5
g/3m2zBljPtt+S5xiWDn9YyJuX4yamFxyXqlsxmkKUFGYTmafRD/iDhst0jgTpHu0bCB+jo/7J4/
HpU9WI8fa1n/V4RDvfWe8LYoXWUkYOdwREdspP4bQk3MB7Y0A7oCOYNohK7qGLvGoHwyto4CjiBt
nu3biTBsNhDeZcH+tP2UL+iDWS+Q59qYPj8jP7QWVROzvWzLvoz6K+ZaNRBkEa2WkirqStduOCLL
UyxmoRd+pUX2O9SMS6MsEPHlUOWYBH5akNXXZoWWnw2gDyOj6XYbtHhLFTVh9PerIfMkioTSaE7J
ek/SGesZsSm/HcgLXDgC3h8wP8YaRJeRYfsUvMhgQV61OUfGPxk3U/6hJtH0VB9VY7OAO7JZiJbP
JJEyd35rXzHrtlvrHmJqh55r9pBKgFBqTqeb8yvYOzqFDVhhHk/w+lH23SKeQ6Y1dF+LVOj2jHlW
vDSsfqX25Hqp2BvE76afuDOl6WD0HI67hOG3VKabz93u0pWhb4ktXzYkVzfKABqLmevgILBMqdKy
43bgk5B1e2AaommnLAYfoZuiP+nFrtNN0PTZjNKphtQpBvi20UyXOj22R54JPBeNinTSNS6Ziu8B
9cETSScRKjlrmGvG9h8SUrPheAOps44IAPbzWVtMgGg5Y9joftFoxfG+xfgR4Pbf1ATGqNjfNplM
0boFlYp8KSNSkXT+UEnJiPb3NoGLinqbqnER/JPZHtI1g6MMmrgMyuU+EDyTOkTTfUVU9RWqTay6
fl1QjKJityCs9YbPKtA9R7uwPOD5c/Z6CqVLWUue9D7Hor2NK3VNDgdxQjFYiszWN2QY8PVsxQ5k
sqV3SjcUrZjsC2Q/mT21YBpITbyXYe37M9UOtsGx1CqzPXSqUHvcRiNf84vuRj/+GVpHuw3QIayP
lr5PzAX/44rH5A/xXYdBruK5BE2d58kkVJiPXO6TvlQI42rbYnve0mBLFET9rCB6SNaBAhFhkXi8
NhKCvtaXbXdJRwFyHk9O5W20GBZesAmKoB/KGRqLYsIOo9CFp3Gkv7zOE8SQYWkkCPi9lUGyk/Ju
1WtnYTyj0BC/oyPbT3w2pGUfhCmpU+AXw+u/ZgbmB2KWtiPH3OBokI8Y34GqeoQjzDM3SkGhTEU5
1aQ5e7iKAfMRQU/vabjg+6IluW4SYEEufbeZaBss/JC6GtguuNTs/VEfOaALUs0EqVgwoRUoBkBf
2K1QZsPf/alm3dZLVY720CBRjxUPQYdZgvaDzRBu0HQwabOmtnlq/Ss533GvNCAmecRaFt3BCXeh
+czU5qnhfJez7RK7olXKQCmJEcALdbRmMBkU1qc+xktSIPIFxXZJumNwaLNZ8T91B0MmevKQ3T/i
i1fjINlimzDb+ZU4eyf6D25VpQJTzA9HL/14OzckGWVm96RHvFTa8UnWgTBxJdB823r5oQ43npGM
ffyRzrmozpOiCBAO/EJwT1hb9RoEOmekmVVIuRLflQKJR6RXxRyLEa5GmouLFimgZZUjVbRWxun9
8EPbPR8VJIktg9CgeDMPvs9YGkhF1TBHSpHo7yX0aVlHzsNovasdi+xqZUYaQBZ2HpmkvX1Gpy+D
VMWBnfKJQao2r/wUD21QQ/7qQbqe4x5/Bltj477avLhpibwZ0Q37uAicuFqJAgepEnhYk2Y7D10j
f4HsXMEfdO+K4Wt2KQfvKlYg8MRdDoFVVr+pHhulc/iM9RI8UB0K2oxqHHlVU/IYf1byMk9XX6yf
ZcWogh9vfOAkGjxWhfPmySLUhO/BzUAgqydv1Dguh28q+E6PCW7Ver8937CC4Hnwvb1bAsMfKC8d
Nytv0Ugb3mb33d89gYjI8vgJA8Q3riHR5JihiRKwrkFlHkUqYPy96JsHpOf3LxRQVAQ4SdBRjaW9
KNvjZVL2q8bM2z03zb84tW4OnUuhispJrJe4a9QF6Xf8h1VJaEJASI9YTgDSWT3YnwzULnfHJpUq
QXMbeXAm0RK3bxmSNrDUbm3VM2zP4k9yJ36K2ply2L5v8rN8/aSUsr3y5HYQyWstpouN0jz0UqM/
a5+0c2F8G5iLO/58kOTIjiw357oCPOYLG0uJFGj5VDTSpEE4SaDh30u9+BzJUosa3gnXHefAz5e5
TSIBtZIuZaX5u0+RqkYWSCiNxq76Fm4AiEfLDqFggSfJ1qyIkAfu7XHZPo7T+VZF9cHAlqtqxXo3
bUiPdwo3up955mXPOUEYle1CyqoIoR/32sAtqSqICNO51oO6RWjUg8sNiW7ftyywQqk5PHeVPqDZ
0C2cB9RDHZDc7BO2ltE/MeRnW842JyzLU18C64TXEqIr0PRVeeTCjGHHpHT5aGH51XpY4G+9/Zf1
TBBhtqwhUPRIhelPPmd8LBi4DnlLBwmGQC3ze2AEJtBKggN5WAvikSzbfBT6alP6NbfBPudy3VUE
vwVsQzzsvEYcpr1A/NQLOJyjnobt5S/h99EGwvlU7/GXrAr1bWZsmvUgD35rUTglV7+eMTsDKAtq
Un/l6h0McNZAE4nzX7h40DLulPZy1l9t0ascyH7y/TL+QmShctPCDagTaFzy6PZ38zmRy0JRTmMK
22eRRKSQFb6ImPDOOFgQlsLNSqkpdUMDUgRomgcuacX4+02sKA+lE9+GJzPyrNTUYDXWj3PvT6Tt
NHerbRUNkg4k70aklriRux0KrDbSwk8ssB8CFWUsgrf6MAdxyj0dd1s0mu41dxDvrzty4zjMR7M4
T3UuvuK5rgESEVizvdn0dQE+v7s3C35w4DPBToeWuZ92a5WHdV8lNxl/ARkhCvudY1kXggX0rS/7
M9C7B+S9ju33kv/Z/7RgHkBVDsjt8NAEFGpqNT0ksU0bIfh5QMrEIeXmeeRb/D7AHGcB6/QE+P8P
CaI8Mm+KaEG7yag2F3gHagAyryxv3zclTxxo1N5tUZWhftKyq/kh6jDcJaRDClITUm4aB+atCBT+
hNUGpwf2NO5XODC28hTVphK9/tYjl0NhuWXtRL3dc/QBcrQ0YRi3aTNHUETvPb0/57CDMUZtF3OJ
dyPhFPPa3AWW9bCK5kO164eRr4I0SbZPl2aATcbBP2jVCFhsvjDEWrDPZ2/9SJSh/q5FKh5HmDk6
tsCvygabIONBd4mlUTi2BMSarlZDoWhYo5G/HHskgZLW6qbaseuOVP3//9dB8KD06atWt2j642st
03cS8+BKp52xdrNpW+dbDSYLnKoo++pzsmIHER9arHE3rJEMuanw5C38R/1rAEOkI5VviNwgeEQU
BH88O/4xnCBCKhgDb89EMgqU1Ly015slMTKLKWL8mVtzZOXYanf6FzfOdTgpylzB5yNmLqoA+1o1
jDhPLJ3Dq5ocbRaZU8bWxsnXvT7m+y1xF6MVfoZBus5rxFe1WAg0WUmIjdDcxUP6RQSw/UGGE1gX
6jwuBsh+qQdWWq6JmH3yz/N6Q+io5uKl/VMJwW3DiW9zkHf/fNY8IL6Cvn6dCotTLEnq7lTNgBBR
1pSa02o87yFPH/dM8fm6Ml6qr6BvinUkP/GNoE96YgxJ2atpRUktJqto+Ifi3ctSJxJguv4oYT4M
8Lu+XlUM/phgzM19E8KvA8Mf9eZsTKe7zx+Y0xuTbGJwOQHdtWRqjCvw/ZOePU7sJfG6i5ankg1o
Kq4DpECCjF3Kz8+oBGbZ4LX9rGiCIFXPrLr3LcGaAPjLNIhlAuZvx9EnbYbielh0Qge4kzNg7KIN
+QjdDOuBo1tacdpMncKG8lpt49qXucNOprg6SQPc8ZSCz+AaGhcLlXtRBan1vcgbGdjR0JyljtjX
vbRZYsxIsihKkwLd3BOeMaOQ4SH2lYwzYXvauWxPQrdgWxV4cKzIjOfQgK9c9fduUsrbZ7uUYNbV
O8jW1mVwsOiS4Y6anFaiOThoSqjODlNjK6GG3Mf6ZV5sRgbzjUcVkCp8pkiUwmRT6Z/A9UYkdjtB
ab+XqCGxbHi8CsSk796h73xnXmtvCNl3fDxIu7aZ7ro5D5fyAzEYWemCm5ErD5/QTpZ/nT+Wh29F
2GOcB7fvliNsKYUlBjkEC73u1q/wPMvdXmKsMuFDtns3P0Ws9nJZqxQ2YD3f4KCneV0nIiDLRZBL
u6TzD7LSE7Ep2c27mOVd1KnBnzMZJWfwvWCrasWhaAWD7MmDHB0NVeWbs+UrtTThDuvcz8UY0OHw
S76kBwdOCwXN5S9BmBifEzZ++9+U5q7/zZysifPCQ+9n5sE/UrftE7RrHfREc9e3BJvFYTLG//Hm
E7HLQ6AS8IqilxTSvYAQk8dSun7F18cTjS91WDeT7dQja61xpfTKb0fl9YyAbe8pgll9T2GzLkKG
nv73u8X2/2m7AwdcRL4phOVNjeaVtZMt5rr8+Ubb9g+p8rPhM1o7O2kOBR+jj8/Qpm4LQdt56O9p
ffWfLrIxuLbwt68zSgsQOZAhdxyog62aXv4vaOzcjl42mklVfFUMdllORkHaJLWXgPweAgcIA6GY
C78Wdd79ojwOTwry2rK1cVLhCuHOO4LxDfYb4pnSaZ5ZmQ2rj/zRVVfrj0FK8skZXhTbfNNLH2ZI
/TIMZzJmuPmwUNCBfiVDte48dnO5EQPlHbP+hRb9ZY6uma5XO8jFgqgrvdPVe1NfZOzDsbrvwj86
gjDCAwSpRCCrvZksi8WXfKkeyoEqjIuxsX5RWk7Xr6MCHqOLqxhwt57oSya2urcPRtxeiCMtaxKf
O789fkJhbu0Rh3d75DVZH91tYuikLxGSTVIYC1hKHu9JwBDsQnWLGJXM4bJHMu3zeS8Hmnqi8uAR
XykMVeyEvhaYSRUD5A/Gm9W9yKzXuvjzZt7drwyDcoHnlUCbGy6gPrtqfOjGO+jKD6KWV+34gGx4
SYzE5BPXxKKhOqsW+tI5K3Y7g0sOT0g3eUTxCiE5etLgXq8mOYhzgHV4lB+eBp6si/MalVGZ4qCs
LrAgBZRLALOtPFZXkexVN6BxvyTrCpdIqbu99CAixL7htWOOOVz3ZJUBk1+pNYNVGfzMztvFItAR
vnZXFpGOpGcvApbiAqw9/u6NFsi2sBZZwYVq4CpBvSPlLTcgYOBdhOJN7yWiwxM+GxK4/3j/7F5b
2+PzVwUKrMNrC1zagRyR9HDscBo7BFLSgqVeAcuuX5aykrQnLo1Fh5igSSpXprCzGDMbC9aI8bkB
8sv8ZD9RByIUUMgmBfVeVXwMfA15zvA2LkyZlYiNt9/D0pptABv1o2YFeZ6vFF9do/lGEX92I3L0
CY22+ek3z6eoVBr3AXL0dN3ajcijVjeQsY9YXz14EMb84NCUHYg/k9XxYvWsQHA+ADzE4m8UH5+L
f0/t57pEEJ5KTjMOv1hzk2hPblv6kJFBvdzdX5heHePsIyzvAVYZ1gvuluf3YwvtDiq2a/7U7R0j
1Zp8M1cvYkt6F+cHhIZIIaFXV1fiCGFVSReQQ7/iyMI1WSoBm+6xntQ/tU9Kym5J9XeJpKHGplcr
c+OHrjLzi/Vjq1+PDxrWQV2xsQSOcLCRyzSdRbFB4fw1MYJDK1J5CTfqk7gvbVUqB1ti8cltZDLd
5qGcPgomLNyq3AY6RVtZQiEcGNDp5gu6QPytp2ftSYQIS9DBNDvGyMhc7aW9jW7SR88qXtMzl6jT
lAXgZB2eq4l4Lgo6Rt1uEc9yHA6L1nAMt6s7fi0lErs+na9sVt4ScfK9KhlxHnENfaN7yQTmc7V/
ROMgBnGJ3l9aEqYDvydivuhkz7K7P3L17zT160I1bolqyRaqpEHKy7JyETDwtsohIu6xk4IGHev+
ykdjZpUj760qtHT4rsAbcEZFsnVS3+R7KjPluylYoUr20vBv8U2RiiiSsiONvLgOamibUNGt1lu7
1YynDgrGz+nZ+98DhTb5rDab3SkBxDGCImqZE2+TEqUAP4qEjGfUyWhHRGl/dvn57bd/4LSiDYZS
OcpMsSCsFnlRXplVoUd7akXfZHADJZb3bmRfxJ1rak9jOUE40XLcZV+UXM59dlMQcFMbAE6wHPWO
eMPdXd3haTXAkz75Nv3phd2mtlF6LUqMcN99kivZbRn7d3uB0HYT/iohlCdAvVaBNuzFr8vY/bEj
a9W83yVrN8CQpzQuXytijaEi7U8VPnXPyvEi917m2iWbF0qKYlEA7bYnWBG96Y45+SyJ+pvV6Kwg
/QYymqKx8GTK5xcgE/QLd9ZeCh9J0Kplg/wmFBVhS0n6kY43uCVuc3M/XVIAEqHum/VN1YmPC29B
mooybl469ugvvdfZNTdrEUjdGI9C1xnOdB7BZBvuJiCICLHm/KxooaFkYeU70+JLJ+CjVYJcZvw+
w+jTzr5IT8Gsq7EyLGMYI10uDLc9hHOu7mxWhBy+QSHvHBoOJ8P3SsdWn2uKvdO3YjcKtE6OJ3rv
piEBWJa1QplmGRqndNtVY2c0PXcp4mQYxjEOcqyKDgqOS/8a8izu5sQ/WN68Z44outMrQ7PewiCX
tirMthM/lKmWH/koK+rRDkOUUja/V4W+xCiTBdzdNY59QELbdHU1n7YGFqXYFvJPVPg9P5vq2ww3
siUCTmlrqme9j/pkTymzd0ZV/s4IsH2k9+/ReyEXlDnP9x6lrYFnnOtlediQAXjE+YOUl7bjWLh6
WBrIs5J9WqLJeakZQPKQ8pbkjKAbkwD2Iob//Y+Qg9AoJl/VnayExBZhpnnUct2wNGmsZ4PlKeyD
CVJ6cY+Q7UHduw7OvrdHr+LvWDiA3x57pDP6Ba98aOHtyCzblIlm7v+ts2q5KHqwfNtGCS79Difi
BC0duQpcOOxfL2FkJnLMUVBjh6jwWBO/4GfD+t1Wtg9UwJkhqgMdlQBJVbBPZ93XqmynNGJhWOto
a7Rr4MtO8O6jGN0V/WZI6b7fnOc8VGTxxaaeZ2ZWhd9vR/JScZ8hljED4ZMe2M5MDUTawEJM80XL
0BNWvJj93VGOa7MFyS2WhKzVvOxxVIVbpdIwj+76mkitjFe5SLxtPYVrJSlU3MxSPZuXcj1AN8Ii
7IVDaLjOJ3bC2NI0qvazQC2FXRgIjotEq2gTJHdfwxfV+edNJU/oVOd4kT0x52OAhMmkztJUE8HO
j2DBretGMqGGlJsn0G7SKgj+0/BcW6R+gMdY034Nc5ucKQ1Lbax3pqaNgSL/bvSWHYGySYfp8ofM
o8+Gf1sTjYEZ6yi2XDnlQywW1DpoUJ+v7q+Ld1EYT5Pw/RzF61ZjftF6IL5j9DCC+WVD6MiaWU3q
R61fTO4/j62X2Vold5hJ/OWSN/UduWGDcbRHvsjcQGeMO+yTmMlgVr8Fo6meESDt5D7mmHKLk5jK
MPaVWc5of6tL/Rkws+73mi7MVMQeHDsNE65hZvq6nkBVRtlnL1FaMgq2yZ8St+A4AZ2vsEKwB9R0
6m+J0eUJBLma/p2B+rFIEf3qwJbghPH30Jrk9iRuZs9wu8KE1ahVOLGvtPCyKthPau+Jk+yTJK+0
bKRwj4TnOM9mo1em2TGiTwd9taTVHqD3PAU5asOYjl+sFMd4sG+kSdX3Z4xf0NXoOa9nD96i2qPz
tycQS/FG9CLM11AQIPQngJHGSMcvweO3OkatbgwhkVG1yh0QNZYwGcxgZhlTcSOKA1NwOaD7LS1K
tGTo2eywVFP6/Tm/1hNnR6RARrPB6Q47VAvI/0r00qzVJJVg9UqGNAq9rYYHPTSesqJTrlZ7X3gY
EwiQpCt6AHGz+9Th848OvSOgOR/DWucLBLqxxcvHYiKv46GiMbRtrEx4eXGI81YIJRWA2b7a9ok5
d2oB0S+wu8hv0uOO8l50rQxbquFGW2962Eg97mtuKsrHTAuApCsgbqKX0crtbm1Pv3WDSbgcFTAx
Umvz+4DMEjMRfvVRygFlG8ZHoFOzqJep6aKwlhfPvlXtiWvs5UPgq/x5US5SR0cEvXmqB0w/pGkp
kVO3PImMVSQI7v5SjBtESmCWdwx58mT88cQrSgC7t/lhIRQsUgZWmOXk2pOcVEQCbuAsnCyLLeYR
mNpxxCgZOJZxG79HbGcwGN/g8D+3PYW3rJW8FWwkj0cOGpgpzWxat1o57aiStjaC6/sCwqkf7dxd
+4Y0M0pG/pVbRr/ebmBNCrttNIq9uoHtDxg9lIH65ylY7LtBtWemfVmAzGXCpv8J2c/ztONpWRsW
pd3cGyljlcr0nWJCtHAeDGZ9GILe/84ysHGvdiMGG0bZzffnTalwqi9qCnXdiaw3QRfgnpEGI2ga
nju6RvtZlrj4KGEjqVakMm4n2bd2tZDqAf46iW3PntnZVJ292oDAZqUe4kQA4uFlJvX/8Ri/Zc7A
ydMJ1Js6Vl98Mu//PIozbRqsCVOYREPFJ2WB8AAn8oKkjbQVQphmHcO6t2Hm/UqMVprhcF1C7bpq
CHzP6Uzpmrth33qEUAQtcBZ6OXbDwgnsZXll4lUi84xMdsJnYDzc8OVszkBhhAIvD8PVk98JkYCj
5aPmxLeiOy6dZhshW7y90Wjo5jKmyqS8B8kKMe+lbwPRp9W+jOIqaO4Nq9najuzOTKyy48shAqc1
+PluKAPs6mnQu/xafmAjyt6spQxgStyPpkoxeInr92V9odCW5rgQz4QORFNyzSrnvJ5NoRQRik5U
QaUxoBisCZ4FOddHa2bmZ5D+FUxyqfnLagAo746l+LJbODdPrfrlQWUPgafzA40jwCqL3YxQ2FjG
5x8RoBWpg2jGraUoQWZfZ3462o15/oQsJoPvsZbJu8uDIQeVxdTBCnuv38S1NQcXozzqQ0c6dzuo
HAXrB60080KfQ4qANZct5K48kfaLa0kwuj3mYFjFfG8trYWRmAzoUpJ5mUUCh3et7L6C8c3x5vSt
4NFpWT9mA3+PX91l3BtThdAjKCPjhzF7I93JGaPOptMAODnLtpsMEpd4fwxI806xipnQrM7kaETX
TyDVvife5pFrb7On3y1pO1ApYqXoQPQ8dSUfwDytFKKzSc2uXIQUzQroP5SGbN0lm9juo7En68Ap
RfbjTok8In/uePDv54EOey/eN1m14JzKuAUW0UDS97CREo3VMkIcjPZDJVWUf+DLW9ikWLEqygWf
SFLPI1J7dD55KmHxRaGXE9haAKOUnXWOyKgsY2Ps6YRxDpNGEhJMO+TUmHAvyeqxjGX0wprDp6Pt
sQn5yJ2Ri8OYjwWV8v4vIrbxDfbqnHt2C2i+RjYQ2UqhqiYTSgUzNWUL2iFcwWUSegP2YRttdE3n
rbJha2lT/+RNoT9tvl9Sk9sMfC5Mg+W2AbeJsSUptGwgflk4e4M95mo2GDaACQk9GDyBkB8rCTY7
Yp+bO3DkRuBis2OzGCs5kMDSax6haVWtYoGx+1uOCJvFG3kbSIDozFAtBUo8Jq8bNtQYPdlkf+5Q
FTngwexfPJabrg+vTNxRQsJye7pttHq2dJb/GbbhFXPaeWNHCNvx1/pmJKZ4vG/bkM4jSPrsylxt
/SAQJl56LNtmZOsoiKMY/e63+BKizcgG9tZvN725fLQq2B2jBObuSzzZB3wVwjvvJQBW2s2enpo3
NSO1F1Oy+HCPcJOq0Q6vI4CcpORO3aBiwS5siFytO0qKw/2fOucFNBR8F7X6P4tmX4kI5czT63xy
iJ5ipkAPDCHgyHbpjmRbJvKlAprNHeK22pQaI3wfLvupt80fnfv+4srpvOxn06/3gFPFGvijFvl8
uyG7dcQ3H4c5yRFB7Gzku7fbdk1C43cCPGZScY7Qv4GqLfO10fqV2a4TvCjRQAOGGSdqzWarhuhR
PbpUfG+HYqLwoiMtrCrSHJTD7qWzT5v2MOk4D5jLBTkpnH0g19HRpbj8RTvMyfzjpHQkSOESZU/j
H1nY1MzQpEL7yec+iRKzbAsSV1UFawUQ7OieQ5MZCAFTb3/J7BBPdv49GzKPsHcRa22gsLXrw/zy
I9Yp9uENZC5QZfcaiq460r2hRNxqYK3qrrnruzAasTRog+6W0C2Y2Nar1fZEkWqnOWfhaU3dxLzF
IbKm1uO9JcHbS0U/dlmjtiQ3+ucoA3UOQtU+GE/gy/rHFvmcd08/jB0OFNJjMw+9s3KVVxLRQIpj
HCuoJToMDa6bpN/dZNSmQfdcjoClnccRhRG+1YoNw4gktSQb0YC8LDfHpm1unJxPuurWBlEuCF+q
pFS1fRmBP55wHj7FBk18pmCCK/Th6V0Oa0IUpXsnwBcYnnDLdr5LWsaehyq+0/uAOYzY8m9/npul
NuRwBWBSpQ3+9scReKP1PnbRT5r41O9zEYtzEEkz1kC2kEstI6DhTID3wAAWuYEQbyzMdicj41WJ
zQpu9CjdUuvtER1PRnCjh/KL0i+3xY8BGk5Fazq0xAOrDg0kviOkmwaE4mojVm315gjPBZWF+Zy/
ALiC5R+SOTkQ6raWGQihny3P87jtEWtUcwMOyU8KzdjnZIex0W7bm2FsYWvz/HkEDz8ZJLB9p6p7
/by1Zz2HS3YWyHv4JlFnt5166isZCZgP0ikTtkWKPID+z5QHgW4e0FnL/QO55666shAfZ+lp09C+
+/clUdS39DvYqtvojomaTbPpd5uQ6YuBZacqgVsYms49RuS9I4zaDq6IGmpdOBeGMd8MV2t+gaDt
i1/IqCDgZ2EwD9vU7wZrz3TDp5NEOeJiA5EXlTn/Lo3rXuDwaiejNVb+eBw6xOPGp6LqyV7fqE7b
4NmTNbytMmTezum5381uyc0VhFQmjJ6ol5BIF9F/lOTqqglSJO+iXqG5wLaW8ta9qcwWZiTFx4e9
waixmSYaGpVAzhnlcKxgLkHw7MGDPRO9g4Q/kFHs9CSOPfiqVPHkhGS+fQsxr1Jo6veYuB6sh5mZ
2im2mTbH9OYsjwQ+6AXU4JeMGyU1IgMNP5ZVgzb/k4Ng4wiNUSYfQ+HetdNdSlaEwCrsq6ohJiT+
x/WJ+B8Y4NNwdFK//ez9PRg3xH2AgTwyRvzOOcsKn5+UAiYum5h7wsUcFLgYk7twODkKY860YrAf
Z83fh5JfaJmQq0WJdAcGmc+HfanTbDkWdLAVBeXmoUptOLipjmlr0eczc2cgpZq8agWVSLTCSstw
2T11TIKAyQRZFv0ohP2NQ+pdF0TfqnvZZQGPTV3E4hAcnpfWTA6l/GWKo52ocZeUGtQNjItc1iZU
j5kEnt45wrV7B+KVPJBgB6hcSfnC1hG0r4R7NG44sApMphoTR0lwuV7MyfIJ9dHY1CqRyod2/isq
LEHw0Wo1KMz3skg2tsf5poGB6WAi+q2VPZEA/4XsBKQotnhbJslXNCHfafBAZycDrx9eoPikwtiJ
Y7FE5RvuzFf+m6l+hXnHegoGq1zVWQP496C5wbuoXBZMwcIX0B6B6q0loLTnRZd0SoMtTriqC+66
vIiU/GeZS78GZJ7j81UI7mToqnvcyjS2FlpAyW3W7olkT2HU1nVJ8as6MKHWV7SOdOC/oPNiS3jL
Jake8wXucClSq07GpQY90SjoVLtA/0kdDW+QCxxAtjGE91jRy9UxwPqVByf98QPuvV7v23bp2a9L
CeltyV2I1+3clbVXSL8lXD22qUjSYvOnhul39Bcxn3g/ADoCVhsUDVOn6rTGABi0s985PmXw0v8s
h346BOiRuMUHYJGBa5ArQ+bJFWh2tpAV7yZOSGsZnqlZvjAWXD8VZ/T0w6cwC7s4UkI0YPkYAJr4
iOODK0mXNUAlnAb7wiJRRrqwqdXTTXewl6a6EYHySxNpUGanr2ZPtKJ4+uXKL+bCqVr6CsE0d7lm
/JyKbcocgUEyuAo+1yJZ4Dp3cMX72o5lsPEIkZz6NwSt/Wuqq16gmiW/ZCxj3+l07D7+SWuZY5tb
TKQ/Tthk9SVgVo58ViuU6EoVKmA5BkEijhosM3m1ac3q5w1f01qvDhS1GLOKaOfrihWS8Sh4RqfM
JoDMtakZY0WCZ03+PzhhTp8S9AP6y+zAGBAF4EwEQrVDw3AyPpW0vrgs2yLKO96Pz8Xy9TSkD0E1
ViPpEhGmesHZDtVvA4KNI+pOhaboIzbjVZiCNVREm5O71IHtElUz+uxOL7rpsuTEgJkoO0D7ksLt
InIS29/WPyQpXDvtR4QuLHs/v//nzbP3i7jQXf2u+AOXs7O97u3NqEI8PrcrPnmqU1X06BBul4ED
o4hF8vWwLceZ0ew3uahCAFkZU1PXAeOy6MnPUPsBWRCBAQgenU18ODFyVAPtIrvb5TjuP6S6Rxqi
WYLXeVBrEY0EyFdU6BawIKWKbJY05yZAvXglWJuGBLOePrL1KgJxTyS05S1jl/YA5zSDgR5qKIpH
ByajbS1LaWE2ejmYKt3b9X7Ag8vB7pRwQpWZ57OoVejUxd9q0VDQpWOGCVg4l6FuTkOwgUM7bQMz
IuFuIoEQ9ooykXCuW2tcBROU51oRigHE8uupN6n9J0rbpaWDNkl+H81eqlCBVQx01sddcQFPLUfu
k1uaFaA/yUiwK++mjRljYj5R1TKgrM5z9KnM+xZQf3+9RBt6RrhGcZEryeWTlMWxINFSQfz4fgAG
pcO/Xltk84oQdvGXsevxEgvc0u+io51ibV5LuYD3w8w7OSHLWJAqO4etUucD5JX/13RtsYsPMie8
Yr1iZwtbvjrYxlXmqqi7KGMlaANrlh0e+s4LkI+DAE1oDNlZxRWlA7hI3Sq26Ansiv8BD8ijBO2X
lcWiuh/0BMppGZMuzZGfteRJcqjksQD8af659peoQdXpgolu13St12U/hh71wgnjR+/HH3YwQCvD
RiJr/0KJrKgGF/m26JLGerdmkWFglB4uiG3u68cV7lL1kB9QfN5Eicq284UtXhtOD8AxGlkkdcku
TLeWG6wGZGzF6rXa38+jSfkM8US77lQASYuA/8dTUDwHYQo++56P3tokZqElp6BNjn3DgnsJN0sO
s2Wpw4BrEWk0PZrd78o/HTtf7gFyjXJ9wq+UfuKvR0DBM4Fs9o5yIjrIUEJx4LMgmJwTNxEBmyN4
uZlVMANKTwZnIzwl2nkvCxQwQBfcoAdLSz0x+2BuMtVPiSjRumThBcwC7kCI0ElSqNEujf7I7cFu
ngnpJH2j23eYHwBwvd2L0o+I0O3HdiwiPoaQ6Gb4BtyG7X0fhGo1xXAloZfj3affBIj/7VaALobm
UwXlm65SAttmGvMhe+U2ZDvBnKHQMcqSrg5Ln2ZWAowwHFeHxhbeun4MjteOGrEj6DDl5a3GJqej
4MoAIyQE68Ds45LutdYhNu3waAnIsv62NuWXWXIu2HJJXuOjsUNUcTCjVhZH5MQhnJrDV5f8lCZZ
YLPmriEMQy1YoTytn13mdjUyY/0+zGrAaY/bwdc/2ScHZvfkgaElLQ7vG3W9XfvGQlWAcZmB6etA
0jmxeRy5X3Roi5Qz7HMoXIJxyouuuBBK3yduHCZHIm7Ksiq9xv7dj3IKEhSMZnDXJIDB4Vahtxhb
P8GXMmSWgWGClBrELOqXKyKQ5pstknecwa/ByRn7K63ZKL9PyzjehsYGRo+i9Py5jLagFav3phsm
a8oyKkdy1Tq76jDoQlMdfJWl+z1CR971ElRCkK+RuWIZ8La+1UqhoG9fiVs52mQIkcqdASmoNKoP
IssIa6SfGkEQBLM/5eLFdGFgxn0kmXFV15e4Y5YlL1CLWVXSpnBvX+huUL0BAJUt2H3BBSflhL43
sTALchFWhm+gLZSQryuENKcARM7dQptBgqG8JMTymCvtP/yBCwAOu+InVcrv3jxVulZnooiQOgcA
+1PX1ZNi5CCOfMnRJNBga44iMCiJ9oLkzQ5iOxzALuK8KeoG8v5NHIdwIGK7beywwfKv0+pJube2
o69wkyQXdtJ7Wdrs81KimauXQvm8bqt2cyWqPMyiizC9DB5kurzXSliQCRhhjbXRRwr61U37Guh8
6DXHv7sQc2zM0PXTUJlPIQIEgZcSxYG+O/WA6J+IIE1NaQowoMr33plFUICR02FZyCoBT17CMk5T
yX+/FcbRAvF9PnO1W5fltdlC7v9XsnVJ0MICZtpZXCI2g7YqQe8jL+7pY7W5f2xGOF1K9JxPSvv3
gOq+AiWbo0QOMwpC26DAkVA8STqMwApW0mdmt49l0FmflhRTZbXLjCYIJ/0XlZRn+a3I8FukmGh6
/FZvK26K60tO4vemHA4PO3sfuJGN+gVfe/KfOIAVsH0J5U238uMc9KhH37zcKa/2e50Cay/fYIiM
culU4GjXt1WpZPsm7oA1v4avg8sPoAJeggtiPXggf9R3FyHiFnfdZWU8CsGjFEY4DGQ5HHuuDxmf
ypaGwOfymCRU2x5CEtLTVhxE2ej9qpj9/fLp3ibl77O8ontU/L3QJbxtyktaFYGwmTFIfRgMu9H+
aB/VWM2t17yUuvsy/BR+hI/Nu5OpHC25hhofjhez0jQDQgv5P5aMJhwlWMJa1Xc2sSbvHP+lmMQ2
NS1nc6PHUc7PXTnNDmh9OfmPBypDH9uVY8J3GOCdy4w658j+jxLVHd0mTQbuhw5lO6ILLwTxkb8q
z+IynSTxlRK/NI6hjdbZmM+S1oYcDADKMH/nYfFxfOTjJbCuSsI38O16JFvAhiiMr6q8bMez9Xhb
MOai0uYg7q49itwFgGT8kMVNFjJiAwO5FVtlhPnA6M1ec3eUo8bLSQaUOHsVMxwWnLboeTSuVuqK
GTdDFjolo/A0MmDJmWOoQJEpJz/EEvellsvZqYR+xYFAJtVFdp+IW2Qtx1GnwALoJjkpLhLlyFSv
D5wY0MCsz9xqUf2Gvu6H7KABAaT1F3R22WXDlKAb3i6kQRqyRp7YLPu8luZwN1FkulR6NJ1X3XlG
BNguUtQGy3Fk00lebxQykoR1S8ImpvCsUic95OORrq9UCTEVhc/YQp5Jv9lEacYYuuFojC20EJkN
jWb4EQN/hvy+Zmdfv0JEYg8QFa+X0zg1vgDFG+xjo4NRJ5WAw1IA4+pxg40BEkUUwoLdGGnqla8n
tj0TX2PqIx0Ge2ec+6OIj5Y9dysBdYTTNsJ9eSaEnoHy9Dp9wCaIQ3MJ//1h60IEfjBLSR/RWnUq
rYcHjEPxbGGZ8G9ab/xXdSggsf/Y8ylGqa5cf1iPMHFA3eU9Q5hgLUuvT9GEyvCKg4rhYuBxYy1J
qIbzYSHDvgTvW6GeOn+iKGXelpDETJrWygM7jUDdrr06cFNb+1+SO85UDvcpQ3B2j1OwVnhP7txC
rtJJpIkGyhEekAS5ZX/T9bVq1KLF3KVPfq12KgtkESqq+VGLcE+byCEUtB2tHt3bwH1OJ0GwbrUD
9DPyQDxUPkWEMaCrfVxhxY/9FeMFY1LfMvINfkgecCyEJlOryH84u3D2+GFFS+xGGylIThEMv0ch
RcfJht40tUqKd4+svmxmeNtLq5rOTDdJxhuTSW10UmwWa6h7fJZlmyEuS6H7tOXO3Bfc51ffoGc+
q9gQ3/sfTFDIZo/0iXns8FirgHY8wTDqO1bHQb23mwqzQJ4wdu6DKc/zBD96ZQw8LxVpp2hjyCjd
6mTDX8y5sqllLKMVyhzeNZcC0A05bJCS6t3zPM1pG0cUCYhz2oDB6gk6YGti1mz6kog3xN1IRqpI
dwjipM3aQ6TV8JnpzWbRaBsjwrhkQxuB3cxvTsnMs/GPCh3ZZeXQ000yam582wxW7ancF6zxL+Ot
A6Ia3QMa9/tY77ovWw4c4pmxOaC+2VzbcYQbifjnrz78RJ8wVUAtIMTf2woecjKgZm7azZ5Kb40S
VSEVk31bWYHzlksAyCHO8MoOTDvUHYoz54OGFoFmJK/m9I/IuBvWT3CRtV8IpcctY+a/AeaQHM4u
u/BK0AZ3LY13WRcrGCooA2I51rEaitq4jsfD13/Nuu/w932n1L0i7Cr9ONRSthQ8JckOIMWw0g0d
4DdylygvPK3rNrdZACa3OgXACaEJlzpwjdLwVgVObiYVtaxN2p2A8U/E9T/lleLIOF0Rw8JHalgC
+55KYuP52UmmSMVrGK3P4m2hGNQB32nH1gLqKmZ9XzVaC96HlCEpGrdejlNg5A5A5yR3bhitvg43
D50nrHHdM7vGWKGZ0WRg1GLDqiaFdf0Tz71dTYYFteki1TZ70846kdoo95JJ1VQeqlqwrrLPGiZb
uWDff0SxW33Xte8m5ylqXIKNnB4WwgGF/l8MHLapYsTkuVdZhTqSbNNYln5UIyMRNKs3zqq7o39w
FOedJXidY+HTQa7OWTCh59b+kpvHkUFJje4/HEh0ja6ucNj1p1X26rwZgKkr6yUF6mYZoWqJt9z0
nGstAoWQ7ja/h9JM12rb2YFx95U+1Q3U/hXT2lfHtnjuWuNqqbLjSZrbjcUQUQA3Imx26Ywp39Q6
O/JWgK4YM3XQuuinCC2pYzAHNqcAQzxunn0zXI0gBKH5zg5kSsCMggbeDESoKkHdJNSGBPNr28y2
ddB5dmdgeM21XV+XLhYqcS5ZQt57H2ym1YJCNBj+WBGokWkmiaWmMkhmlyRimK8p7KulZXz5Em5R
SGbiDkE5ipz/l/Ov8DP86t/wKZFVoldBaVMiDVuRamoBHcpHnNnaSQoFc6qs+uWY8gkZ0NW86+av
oNowZT93CzNLbTl9MWJrW4ZEnJs/CGGI6n6ddXWJ49mm/SG4Hq6cyncIBADqp8LcegwTSLv0MAeX
519N8hXELLL5WHaO4rFFzgq7EXMxLQOMYDsWhXK7gYMmHcNbXIMU194eG1u5ALYwLc+Trk9HPee+
KhfR0YQ1xxM2NknSoV4I0JC6+jJZuWgZw0DCW8HwBfv6zsmlKabspJYybB1DcBa3ui5V8eqn9MFf
IzdrxGfFH6zikcRWur4SON47Lygk3AZBMqMPiZ0wRaQouqdRENbsJKCZAnaMrYdV9GL1ryH7TpfI
Dq6K31Yptsnr10Kh8/iptcSefvBWdGpBgfUU+ws7auFfpgjYRC6bj4KpUUImTV9C0V5G/z0LUs7E
bMNjm0cwTNL7s97dfVKxFcVO5jKavtwoKjiNmR0T/iQFhReq/L1JqJbOaiPyI7CODg0SyBRnHcue
sFYQXCD+kzOmWYapV8/eOxua0wRKAeaw+Ilz+FT+cQZzKUrBqOghdCMHej0wDznRJX9OmyxHI2p1
4tirc++I2O9dxkeYmxLr4cBkufXDHJkF8ZkrF0rU/YXMsDNnuOlw2AgF3UImWlorVzYx+lFGQiSv
qRGYokAO34mplGJGm/OxrcwwvxOAVEozZtvuuE2tD8wiIedTN312snWnk3YZhoaJT2eThlJUyKjU
HEif4+SgNpRHLvL7tzBqCnOioZsMuHUD6C5rPgvf+xtDygxJw40kYYrePJ5i06SqmvHM1jwwa/nv
R89OpFbQWAdlY8q1H5mH0fkO93sdvtXG1V3VLrznbrbIuF3ruwzhJNwJPElF7ODjF9o4OxxDTrsV
VOl8t4jd5bx7YuRroYKX9b1AcBIBGrIdcJVvFFV3MFHbYx23PrMJ1Ks2K5n5coV4VHGt4EUpRaBY
4NiCHGR90RQoavFWMj6w33VkKtLCRwYzzfxfnHRtiA/lTu9b59IswCgGgh4KWPrCrs53vU0s3Nw0
g5TBTkIiNHZCxyqEBxXr0V0Usg1x7c03F05wKSOX6JEEJEfpreg5zsfzjdUrXk4VQa7NjpQRIja+
Ufinohkf5eGVdHQSMhG3bA7Y+qQ/pPz3cGg7ASk8MBlA6NKkqk/lEldWwmbcdjpMCZs8hjoP7imO
J4yWJ38eOZblJgDsYsKBRtRBQ+OsuBnYrIEdPXf2MB7UoD1kON3H6M+wwl5/CbgoUoZaC3v9DpO3
9cF196dF6x27ThAR0sAXDtWyxAP32W7gnzlgypWYbQvNcSiYaZzzB+Qfi1VkukCly/Tr6HFmXicQ
iK/UZbv133tIHZB463pMYXorOvHLp+0iDUIVxSpP5Htux8eFlXwLPCbXndQ5ovTDierqkQKnLvLB
OZa/kdjbkAbMt2ejYPI9LgMnlpTau9a2S+CXCc9J1kEmPKvC+zLVgoKya1X+lKbC5enVggj26pXg
kqoVqXSobmF84WuT2JyTzy9+op7V6N4hezmXiZfWfVJD0CDEVfJ77tM+gPm9fI5nfd90QHowlQ/D
pMpRQXeNDny36MQ5s6bJIQ4hUMGtkLzWWoWaxuqRX2okGycySZUQtmq5Xbfiqt8CwtC6ura2Y0m2
jU0dLTQNrzvxFKBcyGXpNUHT44gitS6jBYA+93KcAInNZrlfPfaL7/raMTrZt3QEwd21QRsoty8v
MIjvTlXGX0gZtO76Uduv2EMqK+O33IFQDLVXUicA7j7d6ZRuLw6pWr/MpsbY+6hlnxY=
`pragma protect end_protected
