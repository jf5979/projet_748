// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:04:25 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
glECd9PYHFt50LO4/XCS2gvbwM+N4w1lzdJTbX2JkU6pnJg1vSqQnUU47B5Snfyl
bZu2qP0tdSsybFReFA1IPa9PuKjk5NJaC/yZPFvhl7fxpDyTMaevoVrclmDZ8O7L
u9BNeJDz1lQqsHV5c23eOYH4bB5ljp3eQMpkRIICP6A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30112)
rAn7ILWFCjrfTKIu/Ev14A9YBpQIWmll7nzI+iNlpx5P2WiUzZJa5tcR9o1k4D44
5y/76dCeUDm4AimV2Qe1d/WZ8nkyryawORvmyfekPP3C0+0jqeEQ8NJC8yAoYhUt
jFFWUgz0uPyXvjl4CZTKBZzKMXiHPNDkYdr0gj77ixJrUm5OyyNQ8EapEyFolN5E
xsXt/D8Fg09FTy+2YOyazg4nJ9RAcVzOdLPRV6ed3L3MVW6fCyTxvDe3niwGrsHS
QvSd+tE0t1kgCFihL4eeZhQt7NdIfU7YrHfjdIC/Q5fsFv5Vox6wejgcx3MfL/ui
VrGtB7Z7OUla1tSVXQWefOpo73bACCf9sTRdlOtxdbyMqk2AeCFLN40XXJLcKO6u
BJmVM4M9D0QFMiQ/Rf0ChVhENCFGbIEGBxF2DSbMNMsqXS18zmFflFuyfVHG1QoE
YV05hcXQuZ/S0uJRQTD0+jgCziVrOZGbg8qtpew+o/9rp0dXecEQbYudxL2U2u0O
w0DGROleM1Jb6GwvRTXgtV0PpQDEHeFWoajM8n2Kkmmd4DWaZ/SyzkKe7U/xU0H/
qQEdTlkFei2bTk/ENkdBg7UaXm46i/PIKL0tQG1bk2f31B68eouxnH0oXngec9ZU
J/nsifIt+l4obTg2SgX4RweIqHHw2lgCTqttvZ2AWVYwmbYrAkV5HDnxNZV8Ny8m
JP+ggFro0JDLKfnLot9unRGBlRa8pU8aQPXgyVDK/gBqDrOOzQtfoSxr+HQxopTW
lWZQqcjhIVevEgHlHxDHTuriDV413AnkpCq66qwxhiaa7q3gqvSHv3Gy6FyWHwNY
WYIaiAfCyYSEQ+uJgO7cjbs0lELtna3YsqmDwi/Qj7Nq7A3R1IEs4l400jppNl9z
vQp5tNroz6oQVsplHAlNO139WgFci2A+tZbzv8dt1Gv1WTr4+U4z6NxFNmsNXTW+
fVxuK0ygBXsHkAiXD8QC+D5wqZ4heXS8F90lotZBGgd44Up98B3Be3/VfTsQ4T1P
X2lFb713qLW9T6Xq+2Irx0C83ZLYvZG3SazAKsqM12kNYtINGMMG05Fej10P84X3
s9dahNE6bTzA1yy4Is2ntWkqEUMk51xYX+zmgpKQGCpTQFKqjAuabqdq9Iu5botJ
P9hJbn706oOocbdRZMdMMmQfxfQSkhVm/80/JzJNFjY9EipnjTgnks8ZJVwHtX18
yjEkBTk6nQ1eA6aNno/B6jLaU4sCKvUMlMi/rBEEZoRXqJ+OHIihsEVE7wCVpmSj
RK7BSkoN4L93c+rvhKg5llqM1NLazqqm5oRSoLWuoBzeGDHsw7gdXcHrd0hjY0f0
0xL2q/5TatpvlCksBe1P+TTPgabc6We4Lm4HNpiRzNuLiUy3ZGy0E/Tk14ca4AJU
d3v1gksD5Z1HbLiaHhr0Pbz4WHcvtJ99N1dytH7S/BmetuhItu3k6TQDy29c5mYo
+JsYyp6k04BtjuRUF1DWulCa+2SSDVKO5YH3LwJxozH14hIUNpfaQNzCq5EelnkD
ubfGfZCXDKnAzBlo1hYlJq5ldCYTlRv/Q8IW7nVUJRDGewqyYb3nbesrhQqO73w7
3hr9uD0oJU01O4JC6bz6TsC3mFrc80An5K3e8T1xdWGjU95xNn+WMmBVrfafgPZf
PYeDd2Omlo7bR5I7Rdt7pKKoLIMJbUYgLZlUr65k7wmvkyFLQz6txpQjvurISRYM
7YGoNVKEArds+QfWRczzPj0nX95Fra+4Eh8Q9sny/7BlNq66mOMQcjweZRoe5usZ
AWwf+p6Fd8HtDeVTq015alXnYZM8jgmLtsiRxH7RHUTU08/4B/MkTUjDsCqd1r8+
Ch8catuFyKECcZLP93J/V8vk71o0qOgZB9oqiPxS7XKOU+u1LoX/TGisAOEzTBad
t2dpwl2isVSezNetdX5Z4R+B52sI+pT1VZIVmanFi6CTpy2NLPLfpnWC+2bOOu+j
Udn1Qnw55994diXFnQdsaE7buE04HKDrXxdLfIJb2ZbzhY/rIavfjv332R3S9MCk
CFS4lErPnN8BK1SAHABUtwH5HF5mV1/dW1z3gLiBL9EyN+Vc/pOqGgyarQAJ19Ux
YS5yBWcc2FqzPR1W0MS1RaHXBA28FTU/0suc6nrOfDmP6fywpmdUkw/xQtxBDRji
hAX/L933qK1ECqE5L1ZM7R83x10CsLT5uLctMCcySMRfdO1fZPQWH70S2ZEgb7gG
AKbKbD7YY581t+HZn5RjCZl9VlajeLyoD3fX5sPU3Au8KEz7+4v/j4irK/sGEbo2
or2c1bE/bVUozVDGdVkEhcosJjWoqxigiz8UQu8zwbg42zSVal1SuyYtyW9VaT5t
mxCRptTd1vC7GqxtxUDYlRU1mbu7Zbt2e4EBmPogEaxK3Hr1+4GUmeufWTZlKYKI
UuBFBzuEDmtiZa40WrEAG7TMPWrZJvaSf0a/nO78a9vnasIwiRa5NQfc2yrEP+At
h+yXRRszEt81S2eQja+LuFM7n1ieQ5vGk4kVeGxNrV2a9ubA233YG69/IV0+9tga
4MBRGg+0D8gUmvyPPWcheIiRhqP3CDfDuHslCDfUTs1xoIXRKsfg7fnb+FG48Hv0
VRSb/od68otdIyHOCzETUYMtSJO5nwyvk6XtRfaVbTcV+oIYt4Yc4CNWnqJDEL7Y
5/DaGwR28Ac0gjUBJxxyJCGwm08TdVcp42RqUMexTIYVh2W+vzaZdDZbFZumbRs/
hCl1aeucOvpO6jylu2x0zk4pWD67y7Tx8A9k7iotnOISH9XnHUlMCXVCBtQD8z5D
QyyxmDPmLcXNKwoTCMw71/oKa+6K6zhUsYR2BZLeR+L19Tv4qw5wGCzVjHsiejkT
7uD2XFaY4KtVDRtjx5xn/mt+AFBs91AtiUuBlSP1ySLOj/dS/yxKp4VctqRPmsY0
28+sj/CA5iinZZnEa3cRP9r8Og/IB9/HnJxw2WWU/tO1hrtVQxdh9bB1SmiApxC8
/vg/o0qy0wIcmq/LsdYgPm8WFYZG+VC6V6goMlODIpA4kc5Jbc7h+d9AG5PQh58k
Y22a2GJoexcS4sjMyZWT3fqAMD80PL8we0lzNZCKP5LHcasVqqYp9a9pqEZkBGKj
Xt7but9kbwyndfcIj0nErEH3nXZls/zUooIrv6Skjp6VeDzuo6+G+9OwXCs/hsTb
N+Cq6C/pB+pmfc+h6hhZwcYpWzX36mrd5oV9EucUBBJu7o5H6hT2tTG54npzsBdm
U01o7ebLzZobPFfUDD5f9loXTOOU/TlcfppbgecfwxspIua8xpYmuQhQNFu+RM4O
I94V6ii/crOmqGC2fRIdEEEiK+zacGBDJsuAKBQEviZW+mz5crXXhFPvDTVzMApt
zsVo8Ld21KSPgpjR3dvKhv+q9KCiCBduUr0FaCKJOdGJ43G3sowMU4aaPB6pLd0j
kiXBJnuUWKNSpIEB5/XdJhISn7bjsTe7LFdhUDNtnCmV4gdDWs5fNwUlH3ost5hQ
xoYAbd7Vdv/gk3kknJVQhju3Md4/IW7q0IjH8LVoK51hWitus7XzIZlUEmuFAqP8
u9A3ostSjRST2chqS4QZ7c0p6xPmbEQONQ4/OeK75pRxhf4T1nB7cKehHNYUvaA9
erLTL3KZOuf1P4vu8+WXH0UF5vYJE5C4amBKpTDqddC2YFGxK3Bfie02kgqfdj3n
UAGIFHQ7qg+uaaqAhHp0KqYSD2B+UUdOPg51t++65WYa5SgQi3AbbmnFKGdXOWFP
si5ylK4qsEkXN7LkwEdBFc2f6e8PMf303ZaIeaK3B+lL7cZGu8H3Hr5YiL8G6IGU
C6tIXuFZo6rqb7VDZHetar/MWb51b9Zuj9CseyEQg/2ods9CYh+qa3R8LVWvlNpQ
vsp3LYt03mY/7IocjxL0WxD8iFoIiDtFEj2FWEqGSqrHZedY9jRzrzpHKhFhqvlS
dCTz8R/PE3bGBHcSf5EMu1xENPVbzA7kJOALIWc3oeOIgNqUJOa86KaRRUbXmFEc
MuNzCsYHSmcC4EP85CjWV7ct2R9c7no2Gs37nu5BwJO5FrtPlGNAeFOBwQyb0qyS
FOALudpWVY5Vlu/D+Mr3Ha5akzyOBsu4StUOxFDyaiwf/rqKDVdQLkL1BqC7OOIu
15sxnyizm9NjboNTZYrvX/f5mltzOQI4wRp7jhWrHpekSSWn3vwmEpAk21+YbqK4
yaC3w4OWOxTlyTFqScgMPb9jkM+AseA4H4iY+5NSJtm2pnU31fwpjXaqiCU0g3nk
Eus+bKzKMwigf6l4N9ArhRSdO2W6W8mDIEIZTOfBoJQiSm8U5XjZsZ65u24T9UgE
2DZJyNT8C0SegHYhZyTxl6w5NUJFJvHu/pTLHJDk16eX3EQrtEXGQSVbLbQ1luZp
G4ye9Pxm5rrydC8DWATqufiEVYIQT/TN/OdxLNIS5tk6IBCd71sPQk4ZihvV0/+E
VgQVVdXrSwtU+oRlkyUA24gpANqFo8ziSGrTzBWAPu5V/8ebjj1UbVupkrGWih+Y
tg9EsrFpUXc+wjpIcWTVhv2e0t9LzxyY4pl6IPNtxcxnXuwEmhu/v98ryfIE3YVs
uhr7QMdJXrRwdH5kVj5XdDsN3ewsUxMnlmojhCKgjZ07jKoeoyuX3BcYJTz1ZZnf
haHp43TL7Xk0dxwvdFrzBOpVR+8NwAqftRm6zgB8PqpOjLnfvRb6D/hQuf9dLLfb
ERlDJjya4SuC6NGdb6m+kRzPFCRawjmGBzH7J5kPN3iI8pQ5/sd5ASbZU/gt3GX1
DRyPYbN6l+ty+O6IL9n5lz6y3UjY4x+gH0bvKq2ufWNQQzo+ui/4IL0uB2Fhe6tA
Pfi9ZX4nXTJG5FBIJlyjdzIszfsLMDcVz3NUp+yjdJZAg7d/2grln8TEtOmAN5Sj
7B2ifYIwUhcM8FPabwJ+1jPlY8ii+rDx2kEZGblWpUogfKGc9SWgI+98s1mSQ0U7
+PZHPsETA5PYLkzxRls9zODnSoNpssPihSIfQdQcl4ie9KrZA4lwCbZzVkGr4f51
C6NasmV9VW6lkmSE+OQ5vKk2jB2wF+YKu3pRb344SPOHOWKBRMZtnRIvP2mGUVPn
HjEZ+GtK0GeMXAIn5k5HINUq9cftkxRzd6JcES5oabKh3ZBYXaDeI8VFw22tXQqe
Kp2YPMm9IH+WUk4gDmrQe6V0JeJLrfpb3YBU8D5XbvPsXujOGScLEz8qHdqr7CBQ
pSfBCE7POzH8TpIwuuQHI/rw3WM9XfrgDnqifG3AYSyx5CQstek5P9q1nhgbh65e
urCYihpjBFE0kCV3ELiB4xo91CwhQsFZBRvBwzc9Sq0B7D8tFRY4veFhS2YTBELA
y9FB+ePOe+cxRIsy2VoK0ivdmPu/Ccfqp7UFuabjX2FlVWqZTX9OezgmsW72rAJz
0svpXEMY+sffiOdbIgsuOFlVmEUr0f4xdoP/UAeHmlBXOUMk/0SKMKuXB7Jntoup
GdvyuZTZBTrWAM1J/JKk7TDZuRQ6dBN4xuHh95DRlh8yklw2BXuZxPOT1fboXgos
RVJ/irlallYKX2hbsfW4EGtIPHDhBCac2dosKD6qKnV6Tjsf9g4Q049TW0pBIC1s
v1TX8+2WBn0riagBgPN/BNd/OYTRVKYg9B8Fx5HzodQzn5NroLdMurNVzr0cC6Wx
6YQB809/C+0w+W5AofXn/Qki/GdZ8CDDY21yFgtLJgigBBvdF0HpTysvjJcLOUUQ
EVwCL8y5eGC7QVViwAWult/c3bbY/zB0wQ9haJk7ZlYxiEU7Tqhqk2vo+AXpJtuF
klGbN0toE6igv4X4/ugVydsDLi21B2kSWfUwzAdEYaTx+bkJD/KkvNWU2yeBGteL
KmuUgHk+lp9FRg87sWshsFj7ttRTIvAxl8KU+wJNaJ+hT/02VAfBHS25xkrdO2+s
oNMwz4FY21x3eaqAA7vIzva5dtW/cxZdrQlokS0gAFJx8K52FapUKne6fHkPuRbZ
iTEPGncLUsbwgBbJY+k8saYArp992ldEzJs65Fhe/05ENapBQAHDaG7b5MJtYHtt
x4dD0hk+cd9U5X/fALHvBKn1kf1MJW7f42DT7RaLUSzWralJfYLpkws24BD/IoxE
qvIoHxjAI8DWiIXI04bJOZnZB6EfIHW7U84rij9QC1Y3JpnWz+rDohD5aQrMSbtO
yKYDWy71SCo6F62v2Zya+ng8/cLnDXichXZceK/YPolN3xN72Kdc3/OXwLw5zNpK
15t+k7HLJIuCXdNxXrLUr5Pdtt3ypA3KjbGksr9LgbO5U40TvsEAA0a9ehNjyXP5
eVoe0bpp874D6DXShaGePUOaDPKr8LhyFLWteY1wPI4KG41uxNzV/0cIUeUyM8U+
ry35ZlER3C6yALaV0Nkkhs1gGu/RDTqA1lOfOXCRt0GikNLKUpNRKm42Sf43C8iH
m6LcdNOi0U0fdvwTnXLpaytRZR6+ywReSa6t6n/82CZBl6CgH9y7wFF89qDXHxR/
xv+Q6sNMxJ6FCesb5/MFqP/gC0GtFfNzg6ek+dSMFyTmeIgearFLfO2vy8kRVVo6
wPFxbPzSCLYBrOmQTxeqtXpElm2uZGW5iqwpl+5Efpd6ZmSLXxI8P5fcM+vb3aTz
c5ob1XRVPtxBS+GRhroRWtpZUOUzah6gnu6Ch1Vw7zGZVS+Od/WMYvN9uXVa3lXF
xbQ/jOuGWrWt6yGEJv4fmbkx2FumtoZP9nIAE45Pv00CitMcXnOkss24f57AzoWB
zAHrVF7jH4FoZv19OgUbYjpK6dpaIr65jUoKNG3P3auFaQlCBXcrwPJiaSor7zFa
pO02V0kUb6M/nKlQbqD6gkIAXzZ8qIKwkrw8OJ/F5jPkA8VqFRg5wuMb5rfSytfs
eQPGY3xVIrCYFHw0G7VVN1+4Eh9kdtQ1WFKvE41m12kerzBg0TSH9fl5c4LdoxLc
feGNEwagMHtc3tkIR3UmTEYUt3EkugaTzaSecEfx6gDJu+izF9320EUsIEtCU8NS
yDUiobWqSjuqJBIphOtqpRl3kb5nUrrkCNZwJt2l88+gbcU7s45JplqXk/jv3wj+
YMrgBoIPf5tTbA3YBmK7drdL9s08oS5aJY4a1JUV/l2NahMviR4OebHqiNck6/oD
5AUwci8eg4aVZtrOPFYZHVLVfGbQT182VagCHWSsXG5Yjx65+G7N1Xpd+eFFItbU
eh9Gi7AUxFKUtU4qC4irBegPA6cgs6JfqNlJT9jfW0UQbGzHrgoJASYtXginHQVW
DQH9lTBTg+Cn92c4d5aJ1Gbj/NTUHgfk2rqWi6Ux9+D3eTPcsDsHyRcEWbtH5s0L
biWuF2LBbyhvLkncONewPgGfVBdEorf7y3DiM//MKNObgcUswX4tsNUE12yfhT5Y
0UYUGge2E+MqWjYeFDrwtJ9SVTJIPjMv9IYoaSlDokcnnNiAjUDXGTlDof8YD+Cr
AcLi3Isxp69/xleVyAGrTlx9bqMbHJLgtCa7+DVXy3NhovRpsL9zSFSd7r5r83yR
rnmq2DmkA6lNxCy4mDvGINMYWVt/ISUYWPJNucsYj8ZVOZeTb9N4MOqu59suGvLw
p05sklCoC2Pg45k3cL1/Ya0q+HhdD3Sxx040lwRe7n7vXIGwqYT7JY6EGM6HAGZQ
8Au0xZWJq++EGSXmI2E+qHWLER7H5Yzz4AWnRsn9dvq1MDu8TFLFqWsoxspdDykt
LXAIzFEcYrwCj0Fw7YijgH9wHv+kq+i6W6WDPFM2TpqPxoGORTcSGAAxuCoX5bhf
uegpteHPmguEvaKSdIrjJgXFaTFdthCSKVt2/rSWEgZddKT+DyOnPbtp9fMiNEZQ
GuwFM8gK3xsdyDwyim0kHqiA6piFJ4th7jt54XPgp5+cs6kllp26dMioiG0+Qkm+
aPMlThH2OQdNSgRLmPuNW4OLqIaYgb5oaTncWSj9ifqneQcSIWjSyQY/S/kBObFR
V+W0B5EjO4SzJmPmgpnc8j4NIRMqBuuyNhVieIosefUkzJjsBoMoEIhorK565dum
8XZ8dlrvFXtQlg5WeR5jvLhthdGEGKPSFAB2XHwwrzHgxPaTtLm0cBXrKa5p9dDV
Pi3Wt24ofyPwaxYE+HBmIMNjBjXSrqqpm7lEN0jfKOAwAT+18xiENaP5EX5hWMpX
PhlLk0Pp2s8YNFJinzpDOX9YpEAP0iUwOEMeR1DjYpPD8ldbuHSq8uL/degv0HlZ
fqgM4C7ZDsYBIK6cZKBVcqOu8P/NaT4NDkVA3IDgMbl6OTLoRcFyiifi4c4f2ypR
H9cBcYgBCbKvtnSKza2liTB9y8++BIABzJNhm3j+3Ww61EL5uMvdpqaumQhNFNYz
Oh4PNGKPOsFDRsNJGwrHWruNKCjWd3y6Dap+3ixT1h5iJ4jJtfISjURc776VHS+5
r48AV7pmf/+q5lw61q+HuY3+2S8xk+JAZQXaiyceEGP7BK7MGVW1X7yKcXnGSOhS
IJyEHBjh8hnoKKsIev4b7h5rdazRclGiB3c4a+DDuBqR/EKSL0c0lRnjz+d6cVW3
+MHjfIvkfBH7YH7PCxmvK5tp5LKAccb7Ta3RLZAbkkX7quiomn3Ry6QhvENxaEtv
g0QyO8tqjjXwft8wyDY+tiyRHCV+mqgYqoPpvWxmIpL7J54KFvsTr3BdWgGEO3qp
jnVmVN+ynFGfhbPO4wx0hEaZDS9VqmADmSBQMDMCzcIc9XWE+tzQYl62xYMToYqe
OkLwKGmpYplxltUCzAANz9ugYZd7FnM05qFDVIogSqj5lcPN76zsE7neSGYbLnXV
rC9SQ118DK6vM3BXmTIINjC1Q4EB210eqV3mCLu1ECAiItRX7/H/te5W7/RtsWGe
Yb/eyJcijdGt0RUWLOlAXSxRHxrtgyDW5czi/mQMNnKUVpfNs/qhePOv7ARxrqg3
Sy3njAnhfpKoGKHoyK13XYEcRaygZFNGDfYG0MYnTFoo3/TXuBApJawn88zpeBhY
EpBCs9rkzgtDSCmQnkN+yXZXqxfZBpK26Srk7JVAX1lFlZlJ4h7MCfhoFSup2WvH
nlsSDge8mfeoVibPbG89PdyuU0h+a5+yWDUWjbniHQFL6g425YbR8fbmt7mjBZJM
7Bl6lhfqkr1cUeDOcf9ohuEui7UsSNyKfsb8OQ5PjPhAzotxvO+0eFXFYQlEiymy
xjsNDGDF++rmd6O5Gm7rc92DjTgcYGrWaS0BwFb8xNigZxBAsjaoR1XhWv5o28TX
FdjDwrkHX/mAt2nwqyEe8EKGyDjsE//Y/3IkcgzN7CbU46ew3gse+FSetJUDa4K0
TdN7DGjx+30mZBd3WPRGNJzmWc6LZAfWr0Y+4fjD/I3QzuKgjDjs7Bgt8TrGslSu
NgH9qIBclzrrDr6zRwq9CmxJD14gLkwObltq+LN4ZqFFHLs2/1k52St4uz5dfI9t
I4UFYJq2v3E9XQvmvVWj6MsH8LiQkioyyXHnznOsYBaBEXEV7VV7Zv4fPoxrslgs
lVplWfuQEGXniIQXgu1Wws3fGvIfw/lDS4HCE4rhV3AZx5X3I7p0tgf6vtMZdBYw
vIdYihiOiyb1byLK6U14eV6oNsdsf4BW+qG4njy1sCUbfCgvaazTsccpo87SAZ4p
CRAums2taqNoKmsoDN21AP4W+HHzOifWGwVBGZLr5j5JFFAMZJ+WPsuc+7KN2/xI
h2j5eZ/pMosYxs+iyFRE5WuiVvuCZVc+UFPsRmkaTUvquzuTNqKkA/NDduuwTiiV
+vk9BMwSFxNpP+qo4Pj6E7vOyt4ti3tDcbJE3PNVzhJnrELMkMeSfE6J1px2sLn/
OJjsDgYaq36i597N8nyDCGNq/hSs0SrlbFNJJBwPVZgFPhIkwTmVRvicdgfhQ6t+
8nEtTTQfc7P25jlz61rBXXeZ2QOOZAjRTYhbJUWwNL32DleJKwBbEVh0vuSxFGzO
LATA4hD4FJNxnAzt0zo75HHPYebNphnZj75CF3uUZSnuwzEXBI8xXrK8jgsd15uw
+f5AX5faAlhJPieYOEoWhceFegMjq5nIRxMcrmBM3gUmbgP2tg6y9JqGRcK8CBBC
sD5769Nz4TuWItz9EPD4oL20LYWma324i4cekkt2gWLuZJhkcn+Ta4CEVMFJZ8sg
EMWXZopL5H03uIIocUfZ9j/RNff8c1dzru1Nd/E8jnp3n+TuzAXguxX26TC36TEp
RfEf4PZ7L6kW5EZWN11UGTk21dLeehmIoeJJPNhKDDJueop0fD7uPrq540v8AmkF
nT7GbWZldIWPv8dEkgPyUeenMbb6lv8BTZREKf66QAUgVBABShlx/sCvjY0qESv+
I4dcbt7AKzvhyGguJ5jEtxajnucIKvmuVazJL2l22JRijPvJ2uuj09Qzx8OaENS+
ONOIQTbSw1Vt1/kniOKR7N45tb6zNXErbIgys+6ileaMskAgSymBt/sc1fHxV6eD
IyWaFzKZ4dxj//yUSuCinSthhFvejg0vi+CJsk2tE1hjJ939E66BQZCZX2UfmnT9
v6f2FsLucVzt260qVKnHPdnG1cjGTk8Nfi1G/tuX5IAYZ3lRmvOwOThn0UO45C4G
QNxMLr8aK7lCyrxvsGUjXWBLict2FYkd0iXEkk49IgMZNOq524g+P57wi/6M+1ie
0Da6vVmLpKKrjHM0H8LHQL96nxTNxV3akYvB8SmECvYZ1Ki9IlEcqBaO1J0MzVni
fB0YAxxHAQreVZYxJdMOa9iOKjr9svMQtoqNKUXV9rznBHOoP9D6S2PcKU7Yksdn
Fgmcd0FbPhchv5WUBny6zfd06v/f2GBzQ6ZPDf26V7hcLHmSYCe1vaObH0xC3OGW
HU653n4vTPKSNhrUWS/3y4IJrjSIs0+b7QV+TL4eA7Z/WBjkQKLSiAd8FjP2Dyv3
VuWCx1zRB+v0Xh29x2/I1XexggkOh5is6x2sLazVyHNURarwLvy4Qk9+j+xSxXc5
n1qq/ZQvrPpGs78NuS6vBGvV+KbNasAsW3s4UWn3cr9oAH1B28niRn1WE0RxzTV/
Y6t/nTrrDYTFGkwKuouNbabBZ4xC7EROrGH3ljs8bhV5l1QX/T7lzDV/nPHRSeRU
tIa2UzB/0BZvQMzhSg4B1CzjRIhitOnesIdx8FixY2wKTuxg1LrT3LT/BCXn6gs9
6q4YIggZldRCsEfDVvUNBpgWA3Gj3ZJmn7qpsA4q6wPHquV94PtF4FEUTh8M2+ek
P8xx2jvoZT6YeuX4CCgISqVBES12mra7VtgXc3wkgfxatke+YFM4oQ9FTnKf6Vue
zL8I+Nov2g2t4rof3fbKSl6jGBTt0hBs7P3Mtk1ukmJL6MPJMsqCipujokqaT8hY
Gpc3U/LYppY7pSGfEJXrFbPVae4Zfnmr783WcqwI7vzCrs0Db+SSSX7UO5/RrbKt
aLwkFEP4LHEejI3nraKLgVHB/8EolDCG2Vtt6jNqEmTDE1gIFj0trOuga/jZm3Wj
0+FpSewtSQ74/sWf4vpqfELHkGiz8ptn+KITMM73J4oKcn6HdJMl+VOT0DWhkYLW
idEWocmR2tW9lNem9SppAPy0pqwOVWVILYMfOgr5lqJ9sS9af4Ymirmd2+s9fNv9
q27iwe7fg8noHNabdnXilBKmrpW/qNI0s4SXWCYDklLKmz3OO23mSp2YhaQLgH+X
PVOHrVxbxp1l093Z5iM5FNkX7oEo0X5RlRuKvhMH632j5Z8beJB0ea8Tr1QciK6P
7kxI/JxmMxY3CFrTrjtMUqfRyL6M91KStnTlhcA9de54Q2pSbPNY+X+o18h99iCI
VQu1Yg3fpafRbILCbUUxwqP83aUIN38uH2ORpCt7vPYQQZw9Lm9CJSih9dZmrjuK
b2/Y4YNlWgT4wopjdn2Kp1WM8l84nRFVI4JRugfY9Xyt5wpNyAwuCsASJyEO74Qg
QRCj3Qyyeo7tfBYDptxv8pbNEwVySHU4yFzDgZEBcPtrwTsceqa58A3vGhaQOl4P
YeDNVdpfXMp1ceBP+EWeUsqnwfr2u1n23DPIjMp3VgKGUWhxj8DAOUKB77HLXL9K
2gb0skD1aR5iAL/OG+ZvFnMeQGe3O89/meAcpvHaWBc4qKDPSKVyGaOiBlO+ohY/
gHMt1voW8ESyKdJFnesUllV30R7AgzKJEio3QiT9kQSon/O/IoJoCGMbWoDpnkIf
iKa3G1S7xXCw35c+YomhXDc63UbArBY+mYON4Let7nZ54jlzxVfhnIWGTVCHomlM
HYlOY7SoIEhsnE0yRrSl/PhFGcC8AwTcgiUbeR9TiSVZYi3oaLap03R01erofiNJ
xanJsGP7snhYzkBUvvIz2W4ur4wph7Sfu5eoD8g0nduEL67TWQUalQYnyWrBwWJA
fiKzue4vIrqeP4moX4awdILjzCpD8bT+wqVeJYqYaESHzPzIp9fJ3qJ/TbVGX80L
m1IwaHWwDEwmEbDovcjIgHU1JTla0h6Aw9BKgKwJjccPiC85k7HHqoBIotMTzlos
4qABdBMdDQSsoKNlSJYh2D2fkieTacmkJofC75RVzS6FHAl3U0c2e+NLoWwhas89
2EQrUcDZUfw04TaN5ebW5UZEF0xuR49i9DmJd464OZXTvAIQPO1FvH+2JxFdT5ug
CjTv5P98+S0AHJ/bjsdKDPcQ3Wqenci9lJz3YZpmlvaUt5PCO+Q+/exrR30jo5fb
j+IaN4L2yppVlnHv8+Q/vEXXkRLujKFS9w+GbcxESUiyzgOFH3VFcggr7FBUudSU
6Y3V19LlKw0b9ducb7HW8YqOx6YE4QA1VhUgoZYdXQzRYQjTzT41c7zw7aZGC+rb
XZM2dP50AkNLqraMfXRYJfgLkKA4KnkupvtZ0xKij27z+wRYPJ4en17N/t0z1uXj
pIcniglj8UFjQFR3/T36ovPXh/o5p72kvOGvQwVYJuYY0qgl1sl+U0JpiHvxurLB
aBX6GCOx0Gdh+2L00f8XpDq/hsun5adZBnPsHrD3qkJ/Ejh2ZPNlfwo/NsHXbkSI
WqcilR1RJ4mprBCdgBOPHc1fBGt68z2y0M7pmi0J8h47JrIdo+AF1QbiW9LW9dKT
+yf+ChXuyylMYaV/q5WWUnwjSAIuK+9j97CtFUoGYBKzCQMddACGtzK30zwHx3FL
rvKBrbksrVH+HGncol70N6zpegQKKr/QMRoyhtjbgsIdfbSmxsY9qwFCn6nGmgJJ
gUKNSbLxXYXPWFD2RtrjM02QQdeKCucCRfgz1oTCh4tpBL09QB4hvYJU5HfpCw21
XKyw5jyyo7hrapOCbzZ3fu5VA1rffH3YJJEBh56yQ3EbsmqYNi3P4k/glko+vL+T
1UvY/a0swlHbj/Ev/Ik+bnk79bG7jXISy4/NGcm+5ynK9vAKr6DsQDuVowMTxwZN
jREct8n4kenqgwHGPbH7CKgo0gJqEYX0xolEmbksKNBPOIIV1x7+NHnU1DiVNWu6
eGFinZytly0ZBorPflMTx3YO/9UiSWQgzFK1tV+8NUL+QI2UyMwcbGINchp1WMXZ
/0Y9qXlmwAcnz3fct6iO9muCOxMl9fl3+yetwQvMB58PWVDuqTXUTpQL5ZqtdH76
+oBPwVTaji4ANvyWxY6/jzzD0JixpdCgjCmGKhv4aXQrw5d5D1u6qPRl76eyKTXu
Zcw4ljZOa5HymXOUZg41S/uvisGWKjd9G+gQMiPOzr+ysL2rUrUS+zg2Hh5pGx5U
jw5Bc7k7AubC8qTCSfXwHG+mCTAkvc++/FqX2jyWFdZeoefhqcw8Yzay8YNZYObY
uSwdVh/X4JSpXu/cnOdbvCXNn7NAtAP9YbFnqS06hsYi5I8CQnfPLGlWmwNfo+Ja
VGnK/VROXEybO4G1cm8t0Aqjs1jlYnrwxP9M/YDaPB5FRwgs2wERCwTNAq/IZqfN
NjNqxadARdUKbhS+gQpugqKkh58Ix3PNxqbbturcZHlGSlx61FzqYmSVUXqPqA4e
IpcSCfUnatRTDaefRvlh1UgfZBPs5hDYGO8lmP6LUf/3AaMUFRtK83b8hrss//4n
KgoGrKVnAchmFvE9WrarRueq33wBZSJ43h0/jNPH9ecJTCvpUjLbjRrFD0jJFycI
HyBJpMba6yg1SumtFkTMGruNB75q5/e/qhmlUwh+/a/FA3PawR5rhXiVzl7ppInN
iDgxkMnv0FMGYJJdanaeaupH7sBo0UaY6vDEtloHvDM0ckZv7FvPT6Kxs4WIcBUx
mTfwC2zf6BgkO5Dz3GoBX83yoQAW4pAzofN9byFmiDav2+w5QiZBHnWtxTP6+hta
FpkbsMBnySbjC+8kZSDchXnGp0CcuPyi/zOnOFeU1J7Q5o0VYr9jkbW8LfQEnzb1
6QIFFJn8YH6ucuybNLmildq6sFZr51eYHuWB1Mpy9QZMyWEcm19NyJOecqBeLgqR
KVwALRDJU4ntYUSiodzxYhtF4XqLUtwf5gb5xGGS0gebEC4GZ3u8Hw1lGNZbNjFw
G/hfI/hoc9CABO8eMvAThJpne1YVRgTCGOEuL9t13bR64cVgNXNpsyivctZQ81qz
n1qcs1fO3jysoRmVTnCxLqfMYzepdxvGgrqdBuexb0GLrzmCGtZC6/c0wj4nrwQN
BgZWuqXLFMQReYywbqDKRW99M/IhkS82eKlFO9VFZmgTQloyAJcAHAM2m9yDtjMP
T78utZN0873Nc1V4WysMx/XE4hC5gzu81CqxEOra+IeWSJ/bjilyutJDQFqdyHpR
OtJmgK94dd6u6OU2TjO3grfkz1+NpfflMi0+5hVd2UTmVKLJB7aG00vPm2/mfLSg
dqcWKZlAvwem0FbUOgGT5Rr7TpIh1NQG59qQekZL98mKWqG/XGpOwUqzSe/VLE7a
MD2ZjwwUz1VTQ3dVGi0t0zZ9ZRV7w2ba1/VDSmLyUyhVnKQpnsSSPG7+w+KZdTAX
TVSrYOqQR9WMZshwuyrz7yWiJB8/+L3yTGMD06+LfXLSeYUCYDVnix/uphdOD5az
PuIqElB2ydzCU7dFbcYY7kYNL2fbRNQDg/F5y4+14+YzaGDdcgiz98dtVTZLqjeU
Wpkh7VfNDe9XAzGcvEH8Kdy2zgXqxy8UR1HQJmJKDUiqPuvdnyDivA8MOfkaWFRx
qM3lMxtSZQWOaaL9cRWYD4yDBbPkjYWIKabW9VtsZFLMKdD48L9PIWcvKy7osWft
yAAXyNdgXWwZS8OyTZLuxgbt8FrKfRi514D5c0NQK1FB8xn/H2AMI5dHe3LwFX/U
SjxnNRBBC0ovRcHlQsj7vsUWX03KNn/3L9sG9xjmGPpVhMIQmh1E/4jBiJFGpgCw
9OxlqqtW6TBIwwX3PNkoeJTC+JSA6qL1JgAhOKdBbeQFa+ZNdy2dauiOy7237F7E
lopV0DYps29CGHyT5uMieofujY7cAjYktuj/H7XqWGjlVJ7Fj2090b2CHpeSl4a2
G3rKVxjVk/X1OsIartHnKKeMqQQJsjjgaYoW5xuSGd5R4MbU2vCmfQXkTyMeEv20
MOGI8+PPBhNpsqgIhjKRace/sjJwxrGZa0py4Jnt5Q0+AK0yKbg2uv+K03GWip8Y
u+PKcjp8BnG6JSzHY0X2glTPIEpNN9uv+ZEcKXVDyE3YDQ23STKkC/2dQAfP+E0X
UGsEc4UO3JvHx49IPhl/aH9Jaf/ExoccXAoXFeIOxMnADvtPlZ4nW6JrRcXcum2V
aR7ty51nTVyGhmpR7t05srRjv5Yt4MIRM1KAk9nM+JSmIIPfyEtfuTxn3ny6Zz2A
go/x43s3482wkG6qjiJC0DahAfSDZNHwTk3Q35wZLGVzXLLIik1HXTLZv4+z7ym4
mYo+BHxtkmBNdjW/DccGGq2a1IvQmu3L9GuAdWuhiazXIYcKiz5bPbPlTRJDUxgx
P4zckCCMeofzvya99dQ/iyYn4MLqJTIXxa3OfHYpIAisi6nPZFq8+HdIN2cng0kJ
0RxHVB3RoH+0yTn6Dozi1VWXop7v7/fJ7jPsx8SLsomjnAIe02cc/3mv9nHzorxf
0OPxikVcp6C1zpNZOw5c/WEbw8yOhfnclWVYfAjSGR09Aow9E04tTugdx/aOxVxV
RGjxGoyrWKIAbaSC1BmojAsOpQ271AGM84qJVekTsrR+t/5+N/jr2Ogp9p6Tw3Tb
fRwUSfiwaZ/BH9Oy89mYkCYYSkI96dL0KKDZLPjIjOm0qhHDWewwfmmOz6WIHsud
Qu704KCVoUkyv2aTgDkG/54KnlxyZ7w5n9CshBFGDezZr91jSuD4z/CH7M+I0NqV
kn9XKF3RhWvEJlWf5eXCf0sW05lvxbC+NRKjAVUarurq+nJbMOP2ngilXL3c9GG6
Mb2OWxZOF+lIpYpk2i3TKbhlXC0YgrMKg5fKfx8OUTPe9Lz+gWLma8RUjQaxuPos
U6tCbJyjewsCQmcTxHDG4VMm8ilLtZqzr1w7rh1XEAUYusG5mI28oA0gmpazrobl
ew2/Bcswib7BfPWzJ5w9pu3obNVUnRoOHf/G2fJDDGLwviuy7lwR6az0Rkye+lPz
Ihgpep6tH/xOCLfvutg0XjhfFB4xl0cpJaPKVf8jrMGhDofgrNk65ZRDpBtQDOJg
4dh1DxqHOsHmNAo/996KRynNlmTT8XHr4thZ7LbSQE7A3QlxIEeUYYz/2H0Eg63N
oE4PifsYUQ7B3PekBMMoitgZcd28y0ibD0w46nNs5K88NDQKHNe6QMX6R5xzzWQs
6jFyhJvOx11Jd7L5VM9EDea1Zv71lDV8zDgImBDcTfpqF/ry9eN97Qx/dILMdKFg
PAT8d2k9uOnfmNrofzCMmS4O4fkuC9okr+8Cr16VqVfBnpvpNkWhaKwnz+6qQFS9
BQ0z2SNAwUn2I81+Srdp4oUGXhf9xKm/UrbuDaa10JUwsmGojwJ3tJn8smkDEMC7
cvwqFbUMNzSPm2fp1xHoSlLJoabubwpbL5j088USypaN30+/Lez7vlRiVgk7r1iC
lNdf2SmL+DwbLh6QQI1J5oPP6YfiX8ogqi+C0IHVQEKbMj7Plf3aE5mU6S2rRcS8
YKY6hFdfjH0Q2XkAyvZyEymEg5kTkT5L2nAIqhd6K+CndjoxSZ2UsafmX6QC2bE0
ut5IeLY4owUuXPWr8NiJqakVNjwizgj2PmpoLZhIWIU7pHBUS26qJwxYImqx14yI
pgAH7KcqSsVvUOZnPD08gJsFsGAfYIUo3SODUhg7/fDMuQovse3FcbUc+DjHDnLg
o7ZzOixdifjc9hbwZqUVrfEWTyiAHu7ASPV1pGJe+XXTJDtdasA4vgyQbeg61XRi
UiCb0EBrslvG6LW7NeZ3/yCltpX3fudw5OwZOaUxlIAsL2AbS22JYdUs0W9NGeST
iGi8y/ODobtlOgiTEV38+L0JTY5IRAOlkuaEYN+bQBtBxgN9om9tgbU8d6UJHvLS
/uBKMbk30bWOzwJ9e+f9LAVp7AFNJB9PlbPy1R02AQq+YiUda/GaG/CpS4QVQj+M
OS+9iG/r0UPNUJDbdREVazzJDUXKXqXlyAjVzV7g+1hODgMP8fZcxeJj2nc+OqIE
LqrY3N1NHXqbv9+x9mv7u+5TJHFMXApCDYMdrD1IBKOsA7erMxosijclrtAe9SWm
ILtQchPGz1RZ4mafILLEqrZData5yx5nn/kcEvCNEW67BUfPe3GUvjRNS6prIRoq
8ou74j/PAqkSydkz31Ma7fzYkl4N+xVVRJtKkHa0nJQKM5Dspw4XU/tQm8ASY6oz
A8HJD5yNQhpBQD6PB/zu12fvogHH9g31ctEHkMfrrl0BLM62xSby4w+a8uMHerGI
RMeEfyvDvEJZernRZDvD6fWJCU9bAqDKdjcrcj67YmECTaQZCjdqAqlNDv6muCwy
KChtAQQFLBOdicNIWqOcyziB0F9hT5jKInUq6KvUMFVinuhecctsAQMVn7HJW4ag
YF6cvtth7nSb1XH4/EVVlzRaktTsM2CgJsg0gNaYI9T2fTv/QJaUUTxVVx2XiUVn
Tw+71USi3kbPgRIDuWiEE5mScOgKHpRqAdvJttyUYPVWgec7iAdHkSf1RMsk+k3D
MUqIUy2nMo5dIsmHBj80McCRt21J2Q5fQbQhJ/2Ha1HkUNYuzoiGINA+YrgTqNHI
Z3VYOv/s0MnLK9aj8Ju9AXxN40/TNad55/Yyx3LjCnco/Ri1OlflL8Rq+laQcLEk
kXc/KmtcaLUzcSZfbZmNh8SxzbNsmBncMZ3kbDcp2MEMrit1OxflYOdJ3EcWv+BF
w78il15sAvOK0g0F+gzMpC5WFp8R9jtELs+X+JY3E45UDIWmytKMPD1dnBc6ebW9
gdEHNVbskkQr4wXr8v9WxUHEhb+x9ZHxxKgkiURBbtvU+yH6a+Ulm2l8R5tM4LUO
AsFVxmRZil8NR2najVHxr8V12blDfLmKB4xgfYcqXWJ/3w7OUuUYjxdUepuCqeoC
S2wDN30NWEYk0IMWtRjUF1E2JNZO4UdE5vWnRUnRqyd9+Hedp43rcv7tCRsfP73X
jsykvwMe31BjbARNKzFLRWiKAYwhloEcPk6Wsizdn2OQLnDCxrq9z1uFFUp9G+Qm
wFHWI+Jxk2nUMBs7/BYHXJ25GplMILzScsu25/dP7VlU07tpgR6MGrrhcc1wugFY
MUNxp7N1vpEoE/K9/+maHZibzPYuLMU3FPfOhI/zskIumE0IBkmDXvMn9A2wnsfO
iZ2AdF76G4TIi07XvK32sTLFxe3NFejvgLRy2aWg9gkLQjijjuo9fWTO5GWW4cPQ
zt1vk5/e/XxwswNe34pyvDPJRWw2bpwMUjLvtWU3Rpi3MKHRC8uT+7vm7jFTK5o/
C+KsIjj5RSM5TVbCdRVajbFSs1wLgYRRZGkBGUY0zAVeTII8uyjcQ7FkWxDBpt1V
L3yMufOMQ63zmY3xK0aiz1GdvXV9a/S1TfSHLkOYTPXGMqEM7I0rv55fWN70bEML
7UTrZICjc32+DtWaqzipdl3hxKa1TzbYF+T4NlGBqaUZGimEfdaxwXGAkYYve1hW
QSt5Ktm280LyOcOBKuX0kEblaCvTbXOnrOaux26S/k8EuV39Gqf/bJ/gtTAxpkCG
EXSHDW4IFoVujDVjT1++wnHGIulbHIFzPUbL02adCZgL8cYfjRYrIetOTxYr7+c5
s0V07pGH16BTITEHMQlWMK1aQS5Blls8ZhaSiL2Z2nZHHps7muxuj25NmRhfxlTi
cq6EeaGrxwVt2ukeOgioDkIKpsh9Gx36/1p0oh76iiXYSATwTK9BDCxZNkP6T38E
DqzuJcy70h3QhzuTqtjGrWQPfOPVXkE8Z6Ut0GhNPIdrFAMkCFHN4sQHL73wA0O9
1l6HwM95+XNX4Z7Ye2QX6plfMg5Nis1KXtt+DbgRTIbsPu8QeSxUpRiYODPr2lbs
JXY+5KfGO4JGBbHFEKrMAgwPTamQLUHKk0E9HIVja9uzVvhn/781W88vszk+M+Oo
P743qtlVvtptn5SoYbrpejXhNiJpd66FfmmoMauDTj7fBxT54HsVlf7GtcbERUlc
A3AWg8/ConGGAcgXYnOwF6a2d8S/3EOWO1GXCGX9GqXCiMqDICrVagmsXT8MSWBW
ubk9JRZkXKvPK619+gd/YcGFw5/WmJukZguci/riQFX+ZN8Di5L7zPAK+gcYrwhm
i4FwtIKZvIIDnabZ0HEOkbt84370FxaTi2fXf+KXVivNiF6kym2XU7M57GgotmOz
qW9RDUGtt0kBi3O23hNppwrGCM4UeEkuKzCiDjJiTAMcuTYUVJRr3QSfb0F61Wiu
v4wQFE0Kal5V+eFW6BNWdp0fMOTSBlOx9ubdl1NWmLt/5iJ3I6/EJ9OYVa6z0bA0
ZJivnOO//5usqRKW7yE/yWdv0XEj+6BGEBCZd9tYNVQeHfMGrS2lhTapplTxK1ko
ooATj7Hrg4KjvFBT8E71ra76Coi4wDuAoHybCzq9TMzn/7JXP0zfSqv7da1pgE6D
MLuH4itr9M1YVFysEuNnS/SFTk8NnCRXo+QeuJ8fUfbIPVO/LGKBC+WnzjUxb5Yb
yVDUh2qLhThk71LOCTHecFBjc0WL32eCcPUprtA/llI4+PLsw+yiDkNm69/bKQKR
rnxRCWMJT8Utte9YrmvzwkHq8uNZQyUr7raif7Au90govVFLrPEFxoBIgBa0F8pa
rqCQt2pgCc5d+ytpQ+xCuN9wWO16+io7dZPpUhkR3fWUPDsvpSYl+/qt/a4lkgl8
Wcnxgs24RK+Cqjapj93tnBBEfRqjs5kTTUu+tkltBZ3ElrPwVuZOyR6nuHE6KYxh
hor45Wdmk/m02wqjZOoNiZZpSWs1Jh/I1aWY9rHDHVpF/m797z0laroBqH5e5iua
UYLF72kNrDPcSUbFkvD3PSQcwzvwvQ1EdFO/WVBdEpO0xj2rtyH5i/buoeSk44dV
fybH/3nibuMpMbD1RRyJpEIS14csSPhY+3sEcXmJtp1y0yq3ALa8Z954diG44nB+
zsCWM3gpXWIR7wSyYzFklW83/38ewDW+qrIB6WXhg+rsPH8iZPOSLCW6aId4bM1e
NlFjrN+0bTtHrjXzwiHUpIeh1KY5DB4dg4L02Uo7ePGq7FSpJ6bpZSQ6zDv6iOjx
An6E3G3wueJT7WkbMp1U8/S+mbpre0MmV7Ud2SxYoKrvIsozncI6ZXMYNY3ofi8N
9fxQSrMjnPypfxPiU4vwbRPHf2JhPRyM28uJKZetgE2f4bmwMcok1RW9vzbLWBQ+
l4S0q4/kMgGGEPFWjYsuDmijT5Ax2gkGzJJfMP3yF9viA6vlnW3VJrmQW7MYq0bw
nSE1NxxOTuBjUXOc4yO3HVIOje1wF1umEXEzg5KritiuCCWFr/lpX6f64oUNxDH8
bPewOy/RjPbo3F+gO2CUyg+oyc4xlPGDnHZPUFdrefjBgQOUfp08fYfB8PpR3VSb
rrr/4e/iOa24TNThKHQ6xT5pL71s2E5hFthGRla9Im5FfVoqKhymuvvLcBdtcBjo
JZ2TbEINZN0HrmhyZ1+zFU2z70BtB7u9ETBtFzZ8cMVJQGF439PxprT5ue0pNKk1
Zs8/JZUvz/82eig7Ox+LifZu95o6wDZnIfAqZGhHk5tfmWDIjn2vFsFgAJFaUG1l
SfX8bze1CIN28Ny/QVjdg6VGLI1q6s7tAfpGHgo0a0JPTmsgUg7vFnu6ecDweINj
lLNghQvPOAjiSF4tePwVF5KRyHT++OPVHguMDdFf9IMEtwl3n7XpMGexQgO5DdAz
KC0zwSndpRNwxnzD1mAQGL73gh6ArvLVAf6KNtg4s7lWhElde4GWdMTpebH2fhsf
IumwdCdx+HmYOXoqYFnHGBEK8iN97883dg0QhARnlQ4n9WYMcJegCY0mLaUVMqSu
7xrpCQoKdD0OnXH3oxt2xBCR0w2ZvE7pzpxgCF0efi5x5Nv/PuliVeOp4bPQsSiq
n/3yS91lXsC+EGPNFf0ogxgYAG610IKJArSncFkJeOFlRUAJLYdu9J+7fCL5uPuq
FPYSddKyVSVKEN3ICDcdGkVXUfL95rYGtBbZmvConN7nO/FspbEvBxTeUvlQEBLP
YQAenEtwZ5RniVbX5CzOGwU5lGcTsJkuHrAkEeDSUFxxp9pPKQAJ3eTOL843uOr/
GC1EUusIU7NVHKFpc6MaWSRAQ0w26N/YMfxeqE3DleckDLfrYj2EuCbMsQc8ulbN
EP8BO1GMB6fKpaUdfYoSMTk2LIJ4bNmyMs1NrY1gYKCKJBy6ZkqQ93PVpyXKDCO/
7t4xIOTLR5rPuQBBJ1XNXzKNeN0nMV6oqJiArYNrE8CTZCm3j6iCSPATsoaXEXLj
NI0BouiJHjjqYYCZoskHsbRprHIlWHbc0QVyjvohI7B7Dtx9MFIP8WyMa37mVgnq
lNK2xBpGrfl6CpTtvHTquZCiMn7DUV+RRUZzoZ1g1KB1o7Gyv1skKaxzcrY3M9ZC
i4FB21hUmGJyWfGsyrPWGALQto0gDq7drbbbp7u5r3NCk3ujh+2mzX/u0RBxwT4/
CUkgwIufmCuOXUaVjp3lKVxDoA9cd5xp4JiaSvv2JmAPKG1OjLlFhwjAQUHs8y7o
S2lUIjsIdO/qsUuG1XWDKxhzWpY4kaoVBxQq26SbN2Vxva7BGnaXrZWowUb0nfgU
MnUAPFzPITNeAu++2Nwq2JElAQIbpQ/ITh8Mzp6Iq1uWButPiQdHH5Uk+scMDaMK
JJ2vO8oaWNI41RzA9Tb4gcQ2LLFBWTdK8p6KVlVBY/0ZIKgJ012S2dfJhZhtxl1N
Ctv5xZ60RkXFuTooNpiZXs0VWWvDKnjAa00vOe7krxxG0ImuBP9+/LGgnd6lUZgE
0oF1pKmu2/zTN9xdGjEVqgU7Y1wT8lD3iF2vxhX6PfLpMWfR2jBVOcDqyg5h7pfb
xkBNOo2vCdNjPsdikYOxAzMAulOt7RMRP0rafo4nBV6JEhmibvygbT+40KUP10ae
IQhyFJthhiGoRexn92dUnleub91Uj4i7sYNwkEOfKHPalMbBUH/Xj0vIwt9Hk+0j
G/EIfG3xna3DaQ2QTvqFi/KpPngpMSBjftFzkbh4zSih/62Htpn61JQocikjZz6e
yNM1tZTLEfATPDlrsS+loZlRpxbptH7VVciFn6asW7UriTRnnSeIAYFkM8xVx7rF
NutiB2ZoFC2UDWbHGesRmlBmj6ckHvelUqXylFqgSlm1q6a7t34as7RUW0Ha6WLY
nmJI4asIFpzHVJtMfnnq91ZCsgAELkSy/XY+Y31ox5dm5X57eqPuSRZgDeM14g55
XonjEz+8u4nAY1QPSB195kMn+y2H3X6MAJUCAjy3PjUlM2hiZ/xHnJYCC9puXfZb
lQLpSKwqBBJI9vl4+b6m1pceRxRwkZWS6wln26rnu4/mkRr8bZuO5Oi851/txjL7
NK+qcUqW95J2AWdbNd0RquCxhHWnnHZNr3H6Z75ejzFl59XGhnWqnVC9q+4YHjB1
ee4OZaHCyvKrHLeB9h6IJdwZxe+qunW24gO9chq4WA3Bk9hQ0eUwXcDUF2DkQ0I0
VLabuCmgyobC2tLFiQ8AGLcF2ystVPi3xRL5FJlBHIjuUpzckqXeU/p6n8pIoX6L
EDR5d93IA7CLUQhJlo8xNUGIAX74C6DXacKYvRwJr9vbaoIQsC5aFKKidjXZvtaq
uU4UVE5q8NkR3Nomxq+i/ubnNORz1TrO6XHwqXY+wqC5+eMNshGnTGyRQi/VyPkJ
KGQF7d/eG8Y8rUbAsJedvByUJ6bP2eqloo222aQ3KrjkW5bx4ONMh/yTR86aenJr
FJdRvTpd4yahNcZeP6wPHGyJqzk5y28BU9CBkMh6IJGFxc6TAU2olmfHcUpo0smG
BeDDMaJoGN/rhuN8DEvq0YOrs71inTHuZWfInQ+qgq8sRT2OvpmQXTml6SUS9dGn
wND7nTjSiB1Zavtx3K1sudSSp8Rm3orz8enWClfD5fDEWEGeuTovks0kajiJlSJc
m3ZWcvZe5GpartTynoNv1MHzwLIbtaGsARvOJJcApX2GXlvv10C2hJKqXJQjAKki
rnzIeAyb6sh5WOenG2NS7TEa/uF84aIVtT/V3uHIu7e+VT3thBveLkCACafhzyDz
uXYrjeGiASkj4UpGZaQFzF9snjLP0VfZc4rrrTuDlgmJRlH7WB9ewijWRlFEpoEp
FgmwqLjpLfxuqAXw/STSO9vgDnNbzPFuBfDRVwfC1l/gQxPk+q4kYmK7OTlFKADZ
eti/i9gKy4kdxjQs5El+BS2+PcuQnYxTnsmDyYggpMh4hd/p1Mfn+ZFuUcvpbVf9
zPUtfObDgDrXaJeQx3+i8fZMMWGxESeli9+sv1JTSp5sAgBjMwDV7oHFkF9BDZ6p
XNkJ9J2Totb2ymorDlkgXlS/c/hF4+e2YEfJbIyxzlkGJVxGpRt2yv1ZxMS1JvUy
dChhVB9mxWCn9rWn/oPas+VPTwB6ovEv6j0sePQqRtz1hxXiYx60oRWUv6ylD7l7
mITEtFpU/jeKSn1opoEwg7Pr0BNH3xUrSxDbSQr0Bad1IFEABqq7GhP1KwRsrCAE
YgYBLjLYj5/xfdTbkbmuhAg6AXzystj78LK8B9hNsTYuhJ3WSQWAMZed5K2YFUNA
vvp6iRehwFtJGdL/pVzId8QBj0hOye1wCGFBr6l0PHegJ65LyMDYWDTWsWzFkF0N
Fv+b+RR1vf1COVTDRo4aeMYE83GXhb7G/rO1xL2xaVtBi8CDaxKfzidsaPNFm37K
OxGx8ZOfvtSjR7klTdaQaj+657yRJypapHhHOXr6ImUPGtXwtpdJfv0VabU8jeko
CH4c5QjiXhdgFCTNrZWY78GwmtgXd3jPr03Ju+bFhLeA0eKTgKtJn4JfeQiIRaYF
m6nR3DiEqojA4DEIY5R17S7dbIse6PeoRQQedF5+JmPWvFR5A1uh0fq8k4ulKpXT
lgNPZAR6vE4FsX8tnCvHJRsMembn0BouWrEjaIrf5/eyj2sshobhC6EQP0G/6+vg
ZOPkxqR+Qy2+AdoG/3TsjFN4l03vkc4MRpfTV6B0bhsZt6qSW5akVFuA3km7RXfJ
uNhs7UOAhYKbCCKyKlWyxfTc1AoNdPWVcHRWz3aJNuJZjW3Qy7dpv75ZSpVcmkAU
UOjpNYXMZYLSEgdb4pg9IYnj6An2gdH62ZTTUP2qQ0OO80QjnI1imqhinWvzk2LG
PVda9q+SABIpMTyr7MQclKK0y7g8Fyr6g5s7OZno41r72ETx5Eli3TVe2YNLR/j6
gAZmpIby6Db9EXFB7sOqyZXUtbgIeuxJAmiP+U9bARAseaEpOmdNgM95EfjOHlDM
4gESY2nXjkBXJpHi71O0VWM8MHSZZmaYV2IyN1dpOIyMqiQ+4I8APXAtAlNXuwD2
TCOtNrOfLnApGROMBMUwGWBbv2wQNH//v/24SNtSwWvuSeOhvNkRsrAZfLoemEsz
4bONLUWpH6GliXHG7pyTAevioCQSkCVpxBPLvoRzegso+ArBJTNDg0xppWxbsBe/
w6LBKpxRiS7N+yhxiogIOZ+O3NWkKPzLKgpnSrtn1CfOj6SUb5JIFRaZqrn8gVDU
QUw5nMAssDLzkjJuqx654RrNXNToSQlxpQTweo42KmO4MIdPVr5nYMuwCSNqYLLa
KhO8eIKdLyMIsxKauZwLEguYjVXOJfs+zLoAaXRZky0DxDuDqx448KB+04CptLWK
qtWMhvTtAxHy6c5e4xuPEOZGvSpnF1kHfTanqzmNB58aRew+uZoxDiG5mZS7I989
+6Q/HMLF7Udbn3rt4u5OuOe0xbuq4lalWZEQuBB6XK9E5lkBKlpLIqNR5JQTzcrx
h8oUauO+NiJeXcvOHY4jkLzhOupmZ356bGTKVuDpW595f9/mdLVQ1s0mWJLg1vaH
LvTJ8p/zQwr0QdDnRMOfMt2YQVlbdp+OpfrYFZUwaB7qRXOlz4AclQAtOmEt4T5E
V/8xkRNXvjrmHGpi35In1kl1Qa2MUwecvIJU4pvr9BDbld6+s9m9iRbpBeq5vcnB
cDv90/+fnm3I4hREx3cL+OXfNvg920gUju5CrIcdXNOUVAvQZeRm2njmcBt5RXWy
tGGEqkAewzAAvHc0zQOKvbHx5u/24g3jKgyckdNNIPa5oMJbWp8KmRQFEUKX3v3m
rbrRbucIwhm+B6pWoY8/nWa7Ptl+fdIx4vKq0pJvt7DKb6Ybgv7n3G21pttZj730
gsLjbwG4XaOre0wrBUuCV6hujxn9RtvbxdJlelkO9TkNJsY8VVv35FL7oQOdKk/m
7BQdraZokzCBBVibd6vViuwI8SVmxFYV6likRsVJI66FvpDGnVUNJnui8WN0bu/w
764VTe+ilAv48Iz0UmgYPZRtsRFVYgyvIe5Se+0j4MWFMy5HYeFKfcjix6gircDa
mV3PvUfb3hvw/tfzqM8xBUiPQY7IdIYAeE08lyFym+/3MWb9BrFKDwaXni6+cqNx
BHUYz0L4NRoJZjsmHgNQoZUkekESlFNT7SeFZWrsE56oh8wNoGlBDIhQVwp7h6VG
MQc/I5nYeuo6szSEGyU42i/wvzKcO/GfvcEC1vT0jblp7s4p4Rn4rofpvXfnCc7J
EoU9b8REbq0SxEjLUs9dwcSb34sSGFcPXs1VXlVi3fcJnk/s4pjr3QMTqlxqmqbW
E3Ur9/4lHKzu0HdGDxM6EbGR5F8hOwIUGs8Qia/QzdFWB8WTBIdWhxiYV6OEObEg
j7lkddBC3RvIG72Hlf2J1MimJeT29eJP4JjXZv9Raw3/5aY3ONE4enYCKFevXD+2
eOYkXbpHu0ef1FVZwGIoLdPEuSibXqb6gck3lByy+j8aSGPpXYJ59obL1W/L62wr
J0c4Gt28x3jr25miBdzVAm6g9c1PQvlQO7Z6oZVmxrdA3eurAuLZDy8S9twXWSXi
uRoliJL+jM0/7Birl0VNPtGH2vsRVFmDJ+fldS3Fh96KU3xYuQuPB9/4OkdMhvWz
uGc/BnRHKo5cFNocoP2Cp4hsJ3E0Bf+h50O6ST0nCSszF5cvBYsggt01HIByo5X6
sNTkjIdd75SVOO0cpVX5x6OMVFdz/HMUinRvdDzcMY0mlX5GUTnzaS/NVy0hry9V
oAuqTjxa60Kktzbb7wAaK7QP89rNW3zk8IbKCkuwz2aNY7yMuJg1WQZCCemupC3g
d+atDGDYIA5cPxKfn5T+62P87ueTe0pWOtD0Z+IRgXrfYHeVfPF2UEJci0meRPVa
r/f4eCDra80xujbTnf19WeTjcoCzkcvBWNSpekgfKSngc1P2zJO+YNZqyi/nE2wH
5w3T5Fe4ohnI0FNHSmbCt7hNOyLb8G3+5P+QrKi6LLZ3pNaSLwZ/thw0mAecOOG1
vz/947TYhwRGDis8uFHLswq3VPhciAAsQe0z4zP17y7Ll4f+LkVdi5umryBin5dz
QDY2bFU2ptGxn3LV5vC+cqrGdjETi2dvbe52eYt6ixzLHcROtnIaVYMriWZpLDo7
I9EtwNQKUsMp6EcMPijl8mDC8V6Nqt7/CRpqu8IkXp1QFoWeYYmx8ixO43Smab8u
r03Iu4Fw6Gdan/PMATpxoT/k3mClhNdb9D9SkJsV76CTv3q6w4o9vehJgSSOT14y
WwIvqBOCcI79V8yvq3yqrJz8JEKDRKw+2fhag6KyaQFGAYPjW/M8CEBibOjq3PsC
E9DQJM4KF8fDyrS2451sIBTQ+eAxsck3LsokGw98IyMcnKHksZZVxCoCB9vUcWLZ
OQMv15pi7gpKmNwTVsPLvqma3d06y5mwGZb2q9EB2SLoU6uzQo9C1CoE+lG95sgR
a+deyhHjtL5gcAorLSvPJT3z0k4OePmayd0jgl8DLz++t/rmJ9TJ1/8HuPihitAh
q8thZZyeR7VL7C4QgMHUVS/L87WsYcklIatEl9tAGbFQSbFxtOEno/Ws3Tq+i891
jqqsIe1PTQveo0vBm8WBlnERfkvEncTUeFanhe30H9+wcqhYz7n1u3u0DGLM5t8Z
u2/I4bY3f8OhiQbHB0BIIzHfegCbYu8Te/GDQiOUDa4QlmHbl7fXtx8S+UG6bHEJ
+7ciK2V1O8cY4WKD2NFoV823TQmOAlIDndC9rHOcSOGHKlvZVgumKlInyeGwgjb6
1HwXGvKMQJe835lHP4V0ujNFeDG/Qh2uDeuKAFcMEpm1G54ZXt3E4FoYB7977XNx
euAAjIOCCti0VGSqeUEqAjLfSf/utk8fqa20DvPnOceF6QPiU3bi4GK+Rc4j5kzt
yg4hD+TA87SRrFAvmL2W2dat+N37WLhM3cL0Dz+GUk5Q2+br+ribqXn9KeRgSHc2
e/fu3h9FnyZ4C/ry8ToFL64kh/59zZ5Wim39iW9HT9XX0ld5TjQNRAnGp2luv1tV
l+DaZXaEvI9R8HGKTzyleJqv1ohmMi7MTs3QhK+s0PhJQ6W0Ywi75YwH7/Q+9loP
klE5rWa3RLxYyn+HhJpYpC2/tKGcaZ69xn4YGv1qVOLGMmU5GyJ56RHM0xK2UBoQ
yPp7rLtZigpi9cDl+EP7JsFJB/lfRhE4iz9Z/C0VGnbWP4X5r5DnWDrFfTJGpHtW
gB2x5g5fgZsoto7kdakbYVwf+pH3DkXuFdhIvLdWH0+VxN49mSBjxBb7G7qBHK8R
o6hYbCyyJGr1Q3JDn2Cace/q4DnZRqYMw/YxblrnQRZqHevFUBTYfKuqz61tvmPG
tZvWd78JwlcNRk5vn4WD/JTq3+KQzXokD5+5FtO6ZFRzN9zF1sjxG7c0C/WKnScT
QIIzGCJIAByEPj2zjexi52AvtTTwCcFRcfXwpEYrprJUHeHmwiDwg2GIKgbMHsr4
WsYETyBrWARMkF68T3FXu7XnC5o2WWFDGPfOiKucJEJ59iFXZ2piHdTuI/HCqHC2
MybTLAQlZuDv07Q1iYZ6ReTKMFhAM4t6Lae+fhRMUUaiCFffzgNAC+uXAH649AwU
/QHAD3kGl2HwQZQ/gpbFCV38/nn4tkTPx65SkiHiL7reBcx5Iwf2QGZqhaVrxyzR
Cne3UG8NvNVoXO7kMitUUYGKtOnqyLAeC3Y1DQUHlTgdgajE/r+UU6tjRsOQOy2c
c7bZkPyv5zq/NfvkFiEoYq3hsP0dTtWc1e+eYjVXMP2NM4sQHEldxc/UJryIje4t
RMrygrVptz0TWr/ulYpHApVUc3XfgncMYE0CNFsz+ieWjq2ooq3KpjTqO2GhSq6y
X+FAJolO2DCm7qKyAKedUoN5sU/Qmnrs/iEFmjipbhI455wMqAqjRjGh/1P/ML6w
ISTk5u5E7a8/9kfzmZaWG7izxVZnOqIjAuFGbrE02WmOtItH9aBGh61GXvnJntGr
J34bY+hnJFhGt0ONZ3+hiTnyivx0LqCmoYdj4Msq+ewIyoDIO1pIdeBxPghxOvhj
6kvLJS7mZyApQXDkhrljBskEID/bdGpmMY18gfK1qRfoUg4A8RVuBLoG3zZtHL2B
E6sD9ogupvdzVbrvzg3uHObQt4E1Afppzt+nejS5Ot2y86fvICPi825v1/a99oQ3
jBH/A+uhTNRAQwBq8z98o5zQROclDoHR87Y8sUAXRdGNzcgwsneALEjs0I9qdXCy
/I27BAaMGvaQv1oi/hqcBbf0yn4UbcfUPsu/vAWMKAZSM/q5xf3msCF4M6vHjY5G
oK9fwIC9K4zprmKkE2m8HatcyzTB/Twn6WtNpCNM0uaAm4ZejtkcZgZaqaTW/QE6
DUZUe1eAY+N/P6sDq1gCKod4smMaxRVgZlPjkCPNtRU+PDRT5lSXn5Rt1Mh7snx7
WvIgOAGYHQPpqblETjzVzrNNEwN6eHHUsCIN5mKu/SPg9d2SpUfunISSzVhpt6Hm
730s5Wp0URBz9Zl0x6RKOEa7mhzNiBCI6FC0hR/i/JA0Nl2AQfmCV61qwR6AvYfg
w8Teb7LkJcA4MsSok+NzE++5HZiS7+fN32yjWC/vba8Uz15MkuEy0r7DvEWJQpEM
ZQJVFtC1rqJrO9cDd/IAchvzgQNalPcO21GtyQ6w0xsSSpwScVdET/oeP7OJWw3A
zcROL7zQmh/5L9B/QUHOaUUrD/PMwU44ANTciy7Ra8DB/Q4Ap9vyOhror4JO0Kwo
joQw6rduRDuh35LN6VyuxThoGCi/O6wKiz9vk8UOc7sMwwP8ZJxCtPpv8TI/Ddfl
b4gvlyfmXTFeiTNGfqRxfI5aoxyB9PuaFPXAnlrEz9+o37RyYdYCZMHxvyJhUq4f
Ipf93P1v4fxbZH6Pr1InhICh5XJmxDxQSQNoJhx2o+Trx9q29nexRNWcxAhGKBh+
PS61JlWpyNvqmiU11XX8MXba8pLhJcFn7Lu4mKibHHZklILHP6eTF1RCw3Swgn+b
9IOmSyhGQ0UYBH7aRpDsj8hTyDdxSBeojN2rhrqOWSFcHFonTPH53aymPPz4gZWd
KyfQQr+/IgJuMKoue+q3cTnQHupInsHjWzkFfTs66mMo9ouztXsaHJxbifqanmDu
2As30HY3EriUt7o3JviSgVv7a/97XlyTxYW0lSJYLuvOH7iZvTgm4z38KmEXTPI0
LrqHImfedKNin5WwNlDfFJhGbEfeVkjEJAJwf89Gav0coZkWYE71W2ZGHBPPXreW
R+cZVdXJkHCc2yWqnC6ZpxcdkufjJyxvXYQFO3Pl/vskUnsZB956vMgtD63nf/px
/xTM52Jo7qPuTYbJB1rVuVDCj1MP3DeP2AyjN/fqtn4IWkNzDebOctZNna1X5PkM
MqWMuVIWZgqKJyFZTXOqPY3EfgLUZXw3glt8FnhpOcBPgBIYk3RtX92lQN6rWG/o
pg4r3CbrD680yzZhnQl/4FZfTYDL2vu+9oLvA3xA4BiyQdWeZHXGr9Se832pNE96
f67RcJ4wLuOUOceWC/wwrnFSEs6HJxuHEk72hjV9yZUtWg1DN9cbAoEgIhwV3ug2
cIjzupsvxlhnQPn8ME9Lc9OT1cYmG2IfhuBLDLU+mzoe85vyBiWpVdARBrUm09u7
hHwdDB5/ixwegSjz+htcfnyKN6qEdr+qDpz7S7jSJbMZG5Ai97AV2nEPWLQl8YYZ
kr6kWDdfoHz5nz21b1A5fKQ3H2UUIYOFWOLCA7XQou4hSbilZKqMkuCAFJZ4cRlJ
88yCzk/5zfQyPp5wwJDacv2mz8QZHz9SI1EDuRpB7r7xASjvE+zsvuMJvO1x/Ksg
knBuK4genaexDEFQL9lbXqn6Mj5j6whzBTrJmajLKzQOkZ0DjYfgmNNARlp3Fc62
OpnC3P6fwJqrPMlw6LcyVeuwcT8w8+az/13e2xBmupI5jrsEeJv8ZYn0M431wnql
Ewl8EqI3dftwJI64yDW2V9zLA5tzGFiys2Eu4JlGVOKXwKrpRnlaqEG7d5P014+J
40pu7WCtqqlLRAyKYgriapZIJOkQv834Ho4uypCxveAzvzMg3wEQxNJdzR1ulKc9
Ntt/V/LFNjJXkAJVzzcHKM9MfbghCaoONORfAbvTD2mmIVeLC+IVDeUL0r3GMHvt
ZeUfTlgJ1bYypEDnPMGZihtsKtK+jAASlS6Y3cKGuvPj6Zt0TWD2qHn8OVR9Dg3s
J+njN/l08qUN70Lx2bSdJgApAnzBYByTicMpGsd7V86nlfcNKnG2fACf/CbkTD/H
YLWAqBNTBEDK5a+2bJt251iRnr9gLP2JN89IvtUR1vPqwBX0j77ZpoPOZPvThLqv
/giRH46dA8RePJIJHJdVD3P4Mhmu7Ypcx5TmhmTNNRcl5EnqRX4H4e8VucxzmN4l
3hNkr+f4a6AneeGp79kEGOwE7SGBzqh9VjrjuvY2gZIkeCVONL7c/WC7QwqUE56e
dcCzfo2l48kGDoRan7zXXradGkPAw12DLgbmYdOmpSSL6AqFSFhzf7x73uqNmplb
rub7N1VneXSrGRml5lsMp96vGa1yuWfQGJ8mczaJcPZOwk7vDxCHabXneDyR+H9X
2+RqSH9DdPNfeXxPXYjxTZutCUHue9NT/YnqPj5tasdsil8rt5cTa4soygY+Q7li
/gDAOc9E9qQH/kLn6BYZld5Xu0hRx/b2KcOPh3GQCm3AmOjqiaFICos5JNi1bwhh
oQ6rjKCchrXG6tfUtjypUAMBz2JsGkKsFHG7nSij5GViTHiHkTn99lHIsyd7OZ+H
VvCBYNoBxXBnRfPebKVmF+aZhfms+90x4agSurQ/eAj8FOmf/1ccBmpy47VWg1OE
svntToDeW07Sn179Vuq/uDyWepndc37e1YXgESbbMNSuYNaaGlGGUi8soBGCDUJo
tJrys9EjYscWMPlQJs82jmjMzAypRTW57yN756egFJg6gDw7r1WBj7RYFJNNh8Qs
TEPGb5k6g7ct57X5LuuX+13X2nZHDqjXTyLidcgQD5X/JVVpd7GTcymgzHBhsxNr
95NoAkzwE1DEbk0JWKTfE+tYcb+X/0FEh40GtZ45KfhF4gsaSLCZM+9F9kWYn7kq
EYFOlWUj+L5/TLFG4hfqxoVO7LDjsq1A0AXKe12Q2q/nr16FJk7uVcpkqJj4xUy0
2ZEZ3CPtFIt87niBykSQW96n4ANCs8uqDqKTVKXXNTUpKRZWQeub5IeQwRwMLhdW
kD8N5h41Um9nGB/6YZ7JuMbpQfKR9AF8mAk4tbjXBsL5CzJsG2le0i8HMxSm58mn
RRhRnHlRTTBdCpujkf8lrWQTgTvIG6wznIhsE4fMDcrpQqOSRFt08ciXQ88bhOJG
YIeMfN24H8bDHh6tDOnEPKhNt+j1fzBxKJUFhpUpQ4Y/T4ha1UOHtoGplM5cIo8L
52kdCPEWDjjdCH2blk8usnmb7ts5ZfszwEHZB4U2uODwHT53mAQFRBxMvTyJ/3Ib
IAREHCyx9zEB+x4ajJWAoz7iQy+LE11BpdVTIow7L/mNBhkU77wLmNlTF1YSyqSs
LLwA53NUoUNVQdjZepZ2j62Xu3ZGXaorVp5UASGNHGiJVSTnGec2dsOBMbcPkRxL
1vIrlMHtOfSd/kIvgu2lXADPB/vVV2EiC5gJYycUAo5rjHFKWRTNtircjLo5kApJ
/qwg4tinNoGUWw+iIQUobf/1fHs9fff5+r+Y6rkmLlTNwpc/3J4H8QkjoI+AVHp9
vYxQyjBCcBe5mwiCnOnPkJFIldXHdOuhhQGJnTZH5Hw53vmH9c7NgayVK3MvuNQv
U+Y6Lw7B+YoABHEJHhail43AbtHYV6zevZlf1s630DKC9njgpVdOdbOOVCtoc8CL
V5fSkY2y7E/pLa4YGWwZbP3+w589LLXakIAWQUE6A4QICeBUWo+t9B7CdQBpmpDd
0iVRSNMT/dz5EzxUBa11vPGMl7jCJaoRDRdL1z4yyLTU11UiGXOnQ9X88I8M/fD3
hi2fPKWgtiXWKlJJUZI01cyRiKe5oAHoIQcaUZta9CC0MhkbM1HxoBCoeFNv3kjC
6s73KLewywZ8F37u0Xr3VzqroMUbVQIkGbWmO74DHzzDDfa7jDmDISKik+DWRUmG
ZXvH9qXWoJNG6O3ZMwvcGgbgLBC9mVHk/ZbcPNCwJqDRQxVntWlLq4CzrdweNEcB
mx9AL57yoTOfZI60hAE1xdhT2ytDEYb+yoaYxzTTderAAOz53gNdiC8s7+AwVV9M
cfLMvP+yYMYkYceWahv94spJeaJcfcScYyFkSrTeb1qtlpvD+EsjYFxAfR8y+MII
uMmyCpZcE6cMRnODku54nQ7kGjsPq0swKaxpPiOSrxEzNUXsKNXlDawLzC/nqrhr
z3eWLnAi7Up4Q9fT87YnUYXiQ3gY/chZhclSNTAleBDKNv5RoTv5kTmHezjiCfLg
friwKRRZyfp5KlHrIV7l7nED6k4znS5MJTCB3+O90e2ZjO6pEtBKp2zqeleW/Z9T
RSBkEnqxBsQQJSj8+ZsUPT4ur+CB5QAwur9VIw0CXTZzc+akqpblbdNBF5uO+EHV
hskIDdP1i+tbuiyXgrbiSBrgJtuPReO1NUYB3d/4Udx9N7V1afe/AeE/GoMJ0tGP
2xPq0bE9AG7Lx4gQGJ/l06DKKhFqbcLMaySo0U3qZXyvu9NiglEVYHqZ+a4S8nTt
Dz5HwNhftl1S8S3Qo94bqzu1oORr++yVSk0RrEczC5YET2usA6cjOaJavm0A2bcL
fi9iRa90Rp8LnEvPCrvl/z4+ZnZdnoFGb6f/TCEKRzf8bEJKLzXHQrsh0JE+WdjP
fGjZHEzorHaIszlqAlk2RQdRH4rCjasmGU2g02zP09I9GjKxX5ngE8QwW3DvVhCo
UFZgTrQJksazS+CXoyhmZ1FlzKE7Ip114cRKD/8+E9Ni5xxUi+RhVeNh8ZJlsKKE
x0WoK0WRBbLc/dROXv/CuIIAtGi1RtH456Al1S9AXzPBQFsZENWzfw9dZeQCFWzS
q7MwRM7dAFr6hnsBPbB8N/hl7wZmoZww7qD7ns8IgwN4T7U3V9tQCOtm8VhoG90p
R2cglI/CPLmGxB21Q/R8QWH13zzYRye8ycldAjaHurg8urVBxougbgBzOlZGarBg
z5pKBqZ8qrrEHH/YdsQanRwvWFIJJQIQNLXwc5TzyfxUSXcnZ76UVzwk17dFSGJL
uFqRqck1DPJNCKA0b4c/u24chDlz6s7IDfQVx5soQT8JbNxECVM7Ab80ok5K0suP
7c0L5O8b/uyvG6Z9UzPxHaJj6AVZ6zbD1qoIrVMU+XIdEXUV8KeH86QdvZLLEJb1
TF61hvrWmw3fhLyTcJaKhRUPFUnvrPThIgnSx+v1dSBCLE3Zc+PxflQfu2rW2nsJ
XVk+OyUUJlMNJZlK4GDQ0ouAVMAdJkjXixFHiovszyPrrYMZG1b3lzGA+K1+j2vH
DrEWxdXhoStX0cde5HqawLVeePWrbrRkyRl9/sjedKdFBX9q7ndkwroBYqhKkQYV
Cwwkk1mUg3L+Y7CA33s5q0vtihQ/uHUGokrv+qCDRaJ108lYsHptEoHsDLl71sXx
5i32Lg9gJehHYzZ9sMCokMLgGZcBnoujd9W5baT605ZMMW7IuyYZkBKTEt/12PFt
ZXsyHX+0bN6I91GZaNasRyNOFcyOjcYDdelu1+v0Vez+y+fxRIbNOId55S6Z+zgv
4Jx7kOQq9dzP8eiB+qUQxCF75cVle6byt5nJCNaYMvPG1jZcAtcE+gll9qwpZcal
PwBnNw27Od2Jn7w+pbujDNQ3SfQnY/hBe4KgLG+OObF/CqrRmy6QJDtiZKD3eEKz
vWOlCXVkuGc4zKd28K1+SD78aGbyesWkGnmUb/m6kYAaLTWXFErwWd0ixahsHldE
szMH7i6DcEli2vJUkoVJiuTuNdm80kbqsA1W/U+lgseUob4nPe7O5v2+R2hCqX86
78FWsQs/yLThJSQ84FJtH8TVXpRUw7KwA0g+C7obdsBuKclbCrQUqrnU7XlXSmvr
S1r3RuZ9ov5LH2JRo2JmO6AqYYQPGnA4L+vILAGU11nGVSfzRMVSzxPz9IRMQehc
EwtM+jn6mQukju5zH+jO6t4uj02v+yIPVKtRKGhvWOI7nWicgwkYpZypGP/t8r02
4BX2UHM2ZwR5LmdDKXaTWl80vPXAgzWNGxyoQlFX2U1o1FyivUdDaim1RBe8a8dC
YRjPWVStCyhqHVIR5dEPPL72oO3KMOX5wzY+Q80LHmwEECXF7MOAKDyCfLUxJ3c4
i5fuJXrH9phtChrjewFx3kXjSJIiMTOZqOP1oYmil0FEJ5M1TEBlaXh8igmBcrY9
Zb9eMNRpBqUZgzN27GEWWJstAn3qooiYj2veuuX99jgUM2saxLKsbS74upWxOYFT
uHU4Q3trj6m8Ng0DUHJuBk/re/pTKk0u0iMI3Jedq5+tF9mCtjZ1ioBALtVyQNHd
hTSiKS9hRfVp+92KgZKrPTe8onibvUVnbbgUhDzXMKEGvdrkvlttYNffAomSTYGk
uhh0TW6ZIbDatZxaxRe4pXCzdHBDJb4VVespgvHGVwssiAWLFBwBTTfmpRghLoOL
FThIOliulIoJg0wBwQFbzu9QEtBVq3AuA2MAc5wUnOsxQO62amn/hJ5AF/T7SAFv
6yKyTurzpjCuo2I9aLrccMBJmLLWzbLfNAEpni48VE5M/QooOJHPo/i67mCemF8X
7dO9eIc54DTDYBAwdRHl5Lmk/dtOJ1NOLXe8Y3JixL0UISolFoDikAkfTyMwKhlx
B0NIQzKJQFD5/GBtJ/sDxWjKKdFCZlRv4VrQ1FXMXCuEep6+IM+L115AKgWjVtxH
Fueu2l+nr6+791umMKCMEsCR8nP+IoN3z5aN5dSKG0NQImRMgIhLGewVHwj19wMi
XJnFvKqiLuZPWXJfdGxLpTk6HR9up7QXAalLoRM/nVN3oYl9ZfogD5oI/X4sKODS
9CNeZlfuCI7En/neZ/fUvJQfU6L3eHYZVKbupUkeyLRw3k6WylHq83FXyhrDiv4I
I+01vcA8ecKoomvZBZWsBd2WHoXzj6jWN25x8QhoGAWazjY6tYef3BLyLdvorO+L
B60t4D7w72AFGP/+yU+8FqRftRw+qbUbb+787ePqSYWc6gqrUsk5zDo+Gv0LoZ5f
EIXeDxYVGMD09d1oFJdhqvQkF75JKt/cfOnlN5MpTxMBb/N/9tCoFxiMrue6c32u
lYU7KJc+odLszOrrvcgs0gg/xXSnX73pJb6r5RckjcHtoNXK/ghRwhR74xEVVmZw
q0scZNd6rgZNjmfet8e7jODsLNiPFNqhPDCJDYaZbKmvu6hOwYCJGupVKk9VnWzs
MekwGXsvYMa9bgiYdX9Yv2GeBD0Jr6AYXxWveNq3fr1K5/VsbNomS7/jA/xBPjrW
N4oERUX6mkg5GI2dEU/6KCaYIs8niL4HeMv8INeM3I2HZwQKNK26SEHRDTUOqd6P
/Wv0grVzxv9vq9zyXLC99PbXJuXQeLxduULYYbAQ6VeOprrTk0uJUb0nYoAugBUQ
O2APEEiSIWLJuX609Zfe5XrFvOBdg/Qzvfw5xWPNDxV09EI9Gf8m+dkYmLicnTG8
fqed6VtRJhPC9SwC14V97upuSV1D6toP/w59CvRJIV78V71q/DiXl69q5bCAbyxw
LmSjDWQ2gVu3mCF6V8mr8XTKIEeUSebMqSzmKNXbPhuodPBFE4/HSAqxWsuOpdGk
YzvZojVZPWPn3K6jOebUfrDXQCWZNMXvNcYto68U32gMDJSL5GrAZXFT5cLsxKhe
LCgc1RZmKukC0uCtWOeJLW2dtFh8U2DYEU5DLeJKP32suZ3DQshAGuyoeb9NM503
eQC/RDSdI+A0jO58T+KuOS74MjS1jHCAeByAP1vknak/iA0gXwpdjLyL8vArQ3Wl
FkdZ6exHOOQsDSBmQVdudiQMtNVOSVZNyXnAt+UMNSgCfIdKCDtrMAPs7eC3T4SX
d7+m6QgDswteUeWMvpz0z7sOGapwCwIqZj6E7zw2oXElG2JI7wXpDPm6VDSyRKVf
vSwLaF/bnrCR4ZUHVjZdwAwDhZemVDJbdE8tDaK0re0rJd42NGxyGzqH+adeHo0/
f66Cvt4zNFjifSxAsNzz/4F1FBtIeAMJMDvhtHPEW7AucXZQN77aqCtPbVUpJWY2
anKkyJSI+H6kXvmo1FIh4bhTJC8XEOOcUVZRUXFEdChwatt5flmIDdCjJ8S6Eo5W
JW0A4huV3Ad7gQ+XYwE0asyJypEtBvE5ViJ7lNrfP8XoR/fuI7YpMSF37BwXTTaU
llRXj6NcT13XRL/mrqJTpxv3ve4pARh1n2+VNrOhRA0I2Ivgkk08OWtgVloAYkEx
2TOhuNvMwg7mTEQmhXEsOCzIIMymkmBVO/kIm3V64Obek6FYY1lO6sTamSUTtMzC
HC/Af7Re8GFiiPM8x26+t4mb1a4s5DtSOGdkvlpvykHIfR2udl4ERxD6Vbx8K/7m
xDrI4AwYspSUmHz/LeeiVJ2ujlc1p57Ut0pS6kvRbt5tupob0H7TwcYedWR3ntl1
2GoK6u/nAsO5lPsIPiMoX2LBvU4H0tECKTdOJuz8shwfkAN5MOP9joMcnM7lkpQ2
KW90fbWCGJt5JMe/c1yyNRIDgwPD+VBMoSVXVxE7GvNkE0JqUgWSbcFpDK2b6RgM
xWl8JNmzHys6ZJnZ5rpgXEgnpWmuxDrboaExom7s24tSMonCmhj/UoHFLqBvIULy
mHcG8z6mjQFRvkvjABTW5veREX7BLs5YqPAzqVgNk+zMAjmOtcbsO3sDzbFmHL2D
l2tyRMiLJpA3ra4COfTr7mCNzl2U5PbgwzhJc1OjzGYM79EAtNJBwt1FeGuRgHpj
+5K9olMzAYedom3FPNtklRVlg3637tXbB8TdfQ7eVunfAx/bOC/w0ZtrV9t/CRAc
JSvSNrTZQml/o7iHgDpUnRulhTjv5pxtpUSrPBGspxsWIw5wLaJYsakYYKaa8s6B
pzOYNaF2krDgMBCzFFvv+p23WGHj4hGeyavsEZ+jZ5k3DfELrh3WWx2GKbU7LX8k
/mRqSeeXh0vvqAilXwYt5os3ng+e3QuAIT7W2qNyKmtMVoc0uCI77ef+BCM8fznt
N840vTWAcF6JOyDnJuDoaaxR77C2srCCiAKaBlnFGP2dghjcE+MS5dvtNWU2CAUP
DTbBbVQaDagsloWWR8WuqLoKZm8r65BHXnMpAmODK+eccKr2usdEUBtGJOiFvQCI
0B02F5h/bvLfI0Eni8YjZC7GPi3WmlAwKG6fu6SaGeFJFgtPVtmCBPB4yVTc8XLL
joM93DImqMdGPDH3/wRnzvs644Gt+6Rb79Yp8rWJ+YPGFsT3s59FJzQOWjO6Qoer
L1PK7oQ/Hwgf9iwf2Ktt+RI89U0EVdq4/2Xun1HFzQvCQJbxk6rcyrT80NB1mN/G
+1VHRUFX01LrmT246ecHw0D1NgoVAuHIT1jLeF09YOsPVMfXmCJrCNb83YartJT/
2dOKccFdkp3LtuuQBAWdfzdNBNIpEx9xb7qbj1KZwb89BFossqVMaPTCyCdg+e2/
3zCiCxC6qlVzQq58Hrz7wQydJyIhIHFHWmJm4QyZvde5nCHFzSx+C45sj4NsXnD3
GRrQG8CCtGQ7yW35DrA9XVtWKf5NW4e49QYmlcu7sKYuX0ag1M4ZmCNFXbkk0h4s
qHv5R+zGMVmKiqE19U52Kq+E3jZyqkvZf1gHvFkE3yE2q4wzyNkJGs1xcFTgBEWz
waW1mrg0YTKndSk7CZ1AbELVVgDNd3UBt34Oa7zsec795fRNifUXtemOqOjU2AYn
eE3cZGakC+NSfkN82kkKEtrR+tFGtyIVfWEYyj2eSJPbjDinXSWmG83zgq+zVqfO
pBupzMqCIOcLiF750jLtJ4sDWE++pjJs+oziu+N+hjPJ0unh4RZGO0NuJkjL0sEj
nft00ecJd6OW5bOJwCXIjC2StuIG4RVRSMZh+rYO2APmxJ5eyd+Ts3zhrbNcmIbq
JStgayVPC2f1P1nzdHALkhGIcfZcBa7ceHPoPH6pHcY0VIrV5iG3C/KDW6WH6rCp
6OLFvGVBxCEsXeLg/StCNmG8Q13a+P9eCUAy2fKVNo2+ndRoaBE960eDSattazfn
AftZu1Jhy0nVzprtYA6pqLPFp2hZzPlURZ/AN9WW7+dZI5OJm0vO8X4Oc/i0eLX+
Y/59Rbl5k8qd705nhzThzAM6X0nliLQh1hex+FTjYdZE6lTgL6yjMXfAt4vtPK7W
KCcA0UI8b9A/F5OdKaI6SSigpBraV7FpstbBBa7JM4ds8Q8gBcbA0BP1EmRhFx9i
7t0dEFcBK2PPYCYSGVLZSoLz/hJYbjAbzE7YsJC2IrY6jb1gsIb3Q9lqXIsqtLYA
ZJxs/ulppsmMTr5fzeJAkHkSEgTL+bov+40pSqv9m8SusBsa5e7P/3UaogVBIQ6J
RN51gQc8AymTS2tLy1w2x+xDTwAnitY4/GBE2XYkjNHyWZz421PKjudqFQD3WBZL
rT6brCzbjyNfdnWe2wx9z5XFNAg4jrDG02Q1tL+Fwdsq/TlaAQXRvzZe4huZjmyO
CdhSPBMPG9pz7QVxA2pGHDbuzVvh0cKnrzTPotDffkYE31AHbDXo+gk4CU9ILA1h
jiOwYSClfFItKV2yxF98rsgyG8PGOFbpN3yUUIAgkhP7a6AqOvnfoKmJr2lNJ0Ho
LEKTL+FsAvPY5SJSdlnjMSqqc3Dt4+A78Lr9vnKzuvNMK9fnkq5Fte5ewuB/mZD8
p+zb05QhZ9UGTIjPZxWDLy7zzEKmLOSLo+agF9RpwVbCf9UG47Uxq2K/l3ncDEIo
WdlPQFhVuz1Nf83TDp2SwO5SGcbKFS06MsWCSGWmpLMJWy58E3IKhgmH6ard/8oD
QqB8hEh2P3v5PGCdNrSYsLf9+MdVmzhJZiIKHP7RSwq9ynO9LOEHsSOXrD0nFlCp
5TVwmG2GIEN6qrQQGgrc5TrC8Z4DS5YAQLMf/JWCA4N46w3P3ssfzPDRlQtrem2s
88ZgtSJRBR/bMWa64DdakdwpqK9Sr0+Ys6lU7hoLt7TImi66g9EpxdNR7INNIuBn
4o2nqGL1MCF6Hz8bdbEycQ==
`pragma protect end_protected
