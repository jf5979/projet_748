// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
wVUQAEwr6flUtbM4Ufawef1hYfYpTLz4bBWrv+F5LppUi8LnOA88k/DGtEoNTublBJkSWuFOp1uE
LO0/OantFRLHH/qVh2R6jnoMMK0OsWi39ulMNwNfWhw1RLTLrImStEJ/ABIkgmkdwYA+90L8t7h0
qsPJf1Z3Bh6rxez96LVnIg2dE5KTVGleCC6TfY+76/thpL0i71EArwbCRPcYwXrzbXkdNFDLFFwG
G7GaJNL0CW0b/IP1MYySdkf+QlUCc9I+q99JcjJiOe6dHegTaXpiStsxrf97I4Ko0brRatb+liFK
CVoyXa5Kg5mfnLKUo1JfJcbTF58TZNU00kypMg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 13760)
TPCJXRC3nD39zvBNjw8g6rIMC4eQJtWFLPuyfUc5XTzklD9ugfBD/jb8kE1YS6bNv+fxSq60c2q8
cqOXBzV+fNnHEvuZa0KtSpFS2Bex1GNKPqbcYsJ6NkFz+78IiVBxjU98nrb0pr9Zj/nR/Od4qh9H
KeWHVcJm1U5xGMZnzPC4RHSG9IIif6WLyD+ybl6udWqXasRS2Df7H0KjH8mK8Z0C6WmeN4GJhURh
bwqikK/ayumKy2O0rkNmXU8Uze53uPTQyrF0rCija5PPlIj/UqW25zHKFyRon+H4CPWTBv7mOC8n
HzMMinLn38jILqormyalK+3HFfJvCofGQYZq0Gxfl+7JPY7fFn6pE+ZFTRY6BOwsN77qISpg8+YQ
XlFQlXbfVHzB2Y1NOaZEtmWCkRAilklawlDt/1isk6JeXruHrqt0EHYU3sFCF7LD5PkWAAlbmdF8
3bVjbZ5N5oi58dXaKaBtejJ3E777FSg7jhCYaKDRdmJOYYrIR66U8Ld3uAGHpBKulOiCVEf9bXRc
eTUJzd1owxK1HaPIwkXgBO/xz6iAXsIUvgSfzWQC9ycrMVWs7bKVQ+1jJ9Btu8P0ZonTfc5hwSO5
Ws7q+oqoJ5otAt79x41Zd0EzsjOrOUb2+LLwZovLB376EUk3XqIS5gsM/rdM4zMMCtKR4ZRcnNfw
n4gVeSYbQ3iLtTTF+3T5UXl6Cvu1zP0fbFV8v4vsVU6UQaA6oMeD/KzZkpdA/h+OQl23uEBSiiHY
tsx68oBFcU9fKFmmDI69YTz9Emkz0nF5OPruP/AlF1uOTQj5/Nd1NlfL0SpwwCTSI+t1JbuSRAYk
FjsXSepV8yjfMROo64mev7GuWRFM+BOJCv8VcByCBGh9FyffMC0jiPy2VU6GTg2omWlW+CqUbR72
4j0E64wYsoo9gLvruB4wxUr/gSGkk43JE1ipzKUT1uiESCWfq7gxL8aYWDL317ZkXiGLbgXYtE3v
4RgGR5XMSACrAQunnV97z65tZ2Qn3kyQZqeOEO9JC/X/JPQt3NTERNNQ0xbOyJL4EyxidckpMv2g
nJvQx2d5xAeGb2/U3YG9sHjFjrMPUVEADM0PIPr+GOdkHpw55ovxTiKsKinzBrWpMveN4ntZ53cl
iyIiibglHEQvG9OrE0eCwcish+xQInao+1jpr3KsBU8ULT5fSMedY/cQxzoV11mpaimqZDf2JRoQ
NCbtSb15nZRLZlnZLqFTWKm18Jysx1n/0TMEnFXTQv22KkHkkDfkmKlYin0ZObV+zBmeO6k8k8Fp
1+LKprInopMLGj1xQa6qysy+3qk8kcUAVemWo0gw+wGZJ2V7EKU0Rit5byisWxXLPsfcVpQnABiT
pLbB9eRQreWxukeWT/x4uKFk63D1oPKgbS/JWneyiCSaWyBY+HKF/Boo7fjQGJVtEYNv/CVusxTW
FvSIc6dXqatRotz+OG/gGydiXbVwX4Y15vEVT9N8fpDCURIzBwNfNvVX+ZyvT0PDfhfyVybqP6hX
GWs/ohU5O+VM8rxHQQXFqreYLEe4pxBN9wmvp2EjAG8Oeah5ImYoRJTJvgQTmpfKmqiXkxRTwisZ
jKlmqM+4LgU8pqrIltkgO5LKJT/S4VS9XWiXF4MJMmV3UEBSA21G3w4HRZP9L5PURV62jfgW18Oq
LWDUqZWK46ZojwyHj0iMlY0suduvM6w1QkCnj8QCPd6CAM6a9HDyiuf0RWAs59sTF9ZuCJuaYM7w
N2e8aO7eoQii7jOAJxFFE5y5e2NW5jmwV6ncLYZr2DDSJi3zZpH1s+oY4QTSnIp+ZCYPd7QwEeLJ
iF2OGtWOLpALVRX3OMoCweYxxW2Jw9/3aivb+HmcScL7H8zmHdUPWzPV2V1pd5J2If6Ocw3VD6Kp
kFADsf9sw/Jv2BRCB2BK4Tqf+vwUGBFxUvzh8t1qK40y/5BwDJeYrMbdK7kDlDB/+WyN2sBUHfsy
DB6O9krLeNVmNsXpRivQUOssJiJsqjxtNLpdDnEWkCBGFVlOtXg1CgFAz1vGOIcYBpTjbD6ucz7t
G3gJVGUevPisQUX33pNzw7lrq0tsdvzyuXLKhEWw/4Zo6ntKttGEfZOGYGLICeCGWz5ghwk5+oS6
vAWtntZ8vIMzd/txH2y+WdeGnLPVFulW0j94BAxaCLmDwni3O/PRpiyOmI9jvclchml9eo+0rwgp
czISGS46WvyXjreXg1Lrs2LA/NIjPNO2qwX1C3TcuFWQB6ATwR+8lwQoZpvzo4BRAypP7yGafxZO
DjJsnA8gZVgUU5X4uV8OT1oQp0eN6aCL8WYUMwIzEDkz1sURyUAiIyZzKqfXZlEvg58wgCLG9GNk
guBooHNVdRyK2R9k29947hx7h1OW7zBiYEfHfq2vTN4agrN9LcFFo/j699uNbRf8U5GNKHVLeo1O
9/jq4gyTx8WrCp7CNgvh6XzU3kFnssz1NjcU39g8D372nrbgv/8BAr74ux5e1p28fwRzyir+Eq0E
+tVwoi1yGD2TpkbOnAiyWIsAoHrDXku719zT4qod/8H8Zp2KsrXePweakPZZ3Q+TTtur1axYhdqZ
SEm+/smbFYIYOglRm+ga091tKfM+t4pagAT1hyM5n9BbOtiESk0YEsltLtvAw6jdVZLdurrzU/aW
qxfyXd9x2npUigjjwn1hg5dak9mTgncyB0M5Jwgpst2vilg9iFz4vTXPbX2spKzHG1/1evB2nNvz
8rdzpbnvT6yMOr59wwnaavY3wl7FU91cYLgihYYgHp1A7jAxEcLe7sEYXG/5F4eDsPX1akV/1pt8
3sRwx7P9ewIBur1gdJWng/eXyueUHKA/Tagu3ynEODSea0hK8TvP6+74xv1i2LT1/PM4+cJk3nDv
iedT5QA3Fx0YIwESnDCQb5g/Wi06oDJN8WJmYQdFz0ELSFJ0MHAH47vu7VyS18J73QQ0GTPXDu9B
soQaaTKTW2SR8umUZdyPHUR7xkIA2+wSxuinzw5DS3NkT+0H7tggbVwCfqzsa46rB2r148HsuCU8
6NIoovP8tz1tx0yqZhvplA1DU2GlA7qvviwqWg7Vspmie8BG71gMZkJe/EnM/pAByoDPJzmx/pre
rzu12FwEKGJk79o/FFbWhFJgkHt3wrytd6SRM1Jrc/x+E7gz3PTICsEScQueRMQBEHgls0jbVk4/
vVSJHe7ZsYTCdoM1863G6qejhz1trXTFIzWrFS6d6IGnKh14tBmtp3wZk0QVnmYwYGVaB1np1LV7
GGPFTBypI1sTGsYo6BBZgi1VXjnnUSVAqfx7fV6X+XY5dQaM841xPs/MOJgtJDjDkAI7q149ki5w
aJSbQleymcjGT+wPrZbGz7O2kDwRe81iBghQnrG9l9gNSDFP/UoRHrTM9q8pU894V96qQxzafB9H
H2jnDXN5KIpMQzxPStWOkTURCWoMfEzX0wGEFu9x5tQbMeHR9+wOfMF/15+O54GOxes3qRPUnb6b
UwrVFZ/J/B1yIfDSjO1ZjOOYVFAuGmwTRocdiXZnaqQuUyf1W+HwofSGiQgZiL02atsnAF+wP75y
lXzmcvQwBdlRnAhKmbq9G+9MEsKHnIJgzzZKWxnBTh45taSWSEyk2pbNXrtmbxBeP0yiLtAFEXA4
VooE0jw9uvtARpYGKMjub9EV1FEoq4/LcwAevYkAldvpo91syUDX0tjxkY/iMQmEq5lKHVpJ0qil
zP/qFsLMhHML8P5HME6czegsZnC0g0Bah0SaxC48ftyRylUykIWrnh4EQ4n0lvzmXSqGMivuVNyQ
dgVDgyLa7oumFCFXNzJIYLFRXdG3LooOj0D+qWvp8no4tHzwd9Q79xk15vXovZt9GfYdFbMGZcXR
MGzR+yzvFWkJOiWomUfo2OQcfGR9yb1nChrT5thjJXgaJ5B//fmNM6RdDkXa7bsamuV//jy0vigG
VdwjqA045xidMf4Arro27NHC1IQRZPElrVXoENGgKj/qKg3STapRzByVX2FHPbUfWZ4MWO5s5t0M
756hBg3kS9GsJ+SN4eayESLMQzXqX0M39KosCwj2kcOhlsLUN4p2XiCK2l9kcsd40SdIGuDi+Bey
K1nkwd2rvLnrH9x6QwmjSzVX+35YfKwQdBhV+tYAb7gsOQTm6WA01gHCxBFwp+bYzVd7XMStm3Uw
fQ7Redop4QrQpeBQOvb96oUPa/XUvvB8Fpcj1T7RNwRtWCboPPy8BQuLufmR6xkK3Xq+uzTK2AhU
Sn6biFWp9eVjltIX+qG+HqzaB9BqEBJr7UCwFZa3ZH+arDCc2X7Y9aFEHOp9wfIj9P0uBrQUUYjc
3OieVMu3qCWAZmJG0AXWJm6CD737oV9R8VhTbjE3zITlAkE+sOP9gzwuB6xgXbuk4/M1KOaHUgA1
Ea7uqn1pGh82YijFm9tyNuUW6TMWm4cVMAmVtg4QQIYJyquwPnPdAuUiRJGpfhujXa/zPqL08E7N
1WV1kyOmGSNNq90AjdM1vzrKpSZktNJbK5niSgUyyVS+j4ipGuuyMf0p/d4b2urCXRErejGQNUGY
aBmUDnytk4EhoMLheOEtrpi1+5FeDnsEemnTSqDwKc/R/3XbM0c6bWjpiAAHjkcqfnkXfgUUhcZS
OaxRQeAO0vWUZd7blHKZO4Kax6iT9vB/XMRBtzMg49L4FQ/8+b2Ep+Zbqy4uV4tjN7qnU1THG9Lk
OGCgO4BDz9WcGaQoc+HYyS4sdxmbyC9uHEXJ/h+8LJ8ms/jC1cxUimCWrUuORVt0vi7EmWXKqach
mQxdOhQNQ/QODmp5e0NIZZNA0HlBpq60/LiosM/BWInDTpNLBIPg5Uj1TNUkrG92I9GpraKMHGVE
dBUV4+IqX5nihEy+7TmK8yeThDPw5Bv+3NDao34QDlY0clGDUCJu3Q+gVnpkIE2Ybrb9G9W7JWuS
ZCryy2XBUz55zZ5Dn7SFDOdqoEnWafMx0C1yOH8lOx2DzS8Mnju4IIWyzbgXCuVJeBlGgSN1Icee
2zC8MD6IyfMtRU0GV8mOAqilY3WDHzqCbr74/tMnTiG7PdkzZ+UKlxvzXeUb3C7Y5OrHA8FSiGFg
W8GUxt6IdHk+nM3cNj0FGY3dCjWJrcT8L1t+WydmGP+rXggIsqrR/bBkwYdZ4uFwkviSIj6+jtJD
URHkTgFPe8dMAjTl65+6kP4RIZufYrxKpBu68J2pm8OLrmX9i0UxwMxM2vv4ahuhmakEpnQfkTQx
AqDkEARmiNZuf7sEzh9Rv4VhVEPWtSvVdjMYyDKpy25IO1eTy+MWX3twWhdEqR0Z0oPnGH7tkyze
FMc3jNECeCjFxeHwmL0ysoe2tzd4jHxJ+npPlvgTiaq9xQgSSELHacSYd/oyY2SS3OgdBVyxDESi
ubk5AVsr588OOuHFFJL/+GHnTKQEQj7tmcGWzKnnxEzMfxuZCVaU1b8m/82iTwndA95CJgMX4Gvg
IqRK6bFsdPdgO1SK4FfwSLZ1VKRAo+akmUixJLP+6wbjJwdD/Y3cNF2Lp4BkfAwk3DwDHuYHzTjS
IP3kGLcEf0D+uDo6UMmIFRnb3psZV+Nf77BDxoSb35StyCbq6Yw/mOcxFXZIzzwaK+jxBrrMJQhy
0tFFIGhPbv5jfTYzLsTke+VrhntKp9fEQRjpkwsH6GHI3Dg0mdZ+JMvhXfhuhkvTGK1esHokWzht
7isQe/2Ea9uQM2uY+cgeAG+qTizYRI5E3Fg/wtu5R/FMvLQpdIjziTmY05RYNHyHSebRU9hinBNW
nJqfO0gL7bAtt1gG03NdqJ2M9QifLV4JPiMLdQ0+ohFH9wnsrekR3JIOPuPRHj31zHhCDNNEsSJy
Drith49M5xyT7MqQ6YIj7akYs53UzuS6njucQiJMn27L0L3px5CRmaOmKqhNwmL3RZS6zVy2En0B
33qCcBrNKtEN1UlkzNKqvE3AMfZYeyFt4b0JaEoyVQMnMljIZnAku/9cCGzUFbas4s3yHJnpxgRb
yC5PNnjgv3mTjlWrpc4VSe8WkAQNoXM1P8Yj7eTq3CcgcNIYDvWmic+XiAyxEOE9+LBq+07xAIGB
Rp3Y539+GSgo+XUliwYw5DAoNRZtbPBbdzbc14kjht+VwtJUO4mh5LPAmiPt3Jf6QCKndX6a4s7q
kF3NjKtB/RJe5sEGjt/f5m+R2rwK/aOzNoiIpV0QIOEaN1bs36wQefRa4Jywnkb/fDVbwCZYbgYq
r0Ls4Dl105mTbd+PFlbDqwuJ30niRBCVRJ1PDCBvcGzffOe/nTxOGTSHtWFe75QIRM/Ahh2sgccI
OEu0yh7d5YZRhHfRm2ZorUe8uqpWy+RE4IRHBnUQppew4vCwDM07iiKTY7y126EnQg9Xs5gHvtZq
sncuSAaI7t+olx6AOOZyF4ft8ySxarpHjLM2DCAQDXueR3eDaR9HXjAL6SxrrKJ0tYYP2KPbSFdD
MQDjtGrbsia4rk9jjejSLHx1F9W1caa1UbonQiXNOJTQUJCTwRZTVBwPBdOTaP9ufU9yzgqjjt5M
T6rkksa4cRX9zYrmi0WKH8sN208OxhYrHZ6aQYY6EhlCOWwHUWfavJ424ry3uXdMtxnpjp9ysEoB
4PGFCCBbLBXhTQoKEl6XZIxZsIcr0zds9gdZ2Vi/vBHpVlRtq3XoJ1Q/5WI+00ncXK/biwVBemuJ
hjcaHZ5FNYMZDkmilGWTvgVJWoX4CUF34Bf+TJGoeuJorO0CiBuGiyvJIeYVHWMVaKOv40T8EGNT
IkP99gjqk0+9lDMBHIX8zfdaMs/5Gmkec5NoUvyPv6wfm0xXjnmEIIgxMmr7i+UIJIkdGuuruzm3
7PMr7e7NMxR+gWWjXc/62YcILnnzgjRdkiInfsLhh1sj5SrXyI2V2Wg1GKrQNT5BdT1nCjSc3MLl
Xx1ssYqr/bZZXqhMJ7hueNtgJhd+N/w7jNawraaLBJ2Hqy8wSuV9Qoox9SY+cb9G2EVOy9ktU5LY
Sb+SOVvqkMxnD9BW0eDxDKjlHSTpgDODM9XNY/ZLYD1c1IY1jdOEfnORZGuO3GYdH6f/2hFn6M+Y
kM9kDB+0XboXMhNZ9NqgI5Jt7aH8xPEKfdaqURTjRZtivBRhR3NrRacf2RkVd/sgA7GR0aUsYTWq
8nUj+q++ZS1/SO4vgQLFMasShf1MWAzNlvTmmnv5zPXczlDh+p2lYHh1JXiwbfHdP+FrwgITItlZ
yvmagOuD4/YZse6YJ1ydMlIM+bnWs3y78bCrB2OH3Pg2kpLkEOyIkMsE1NB6Zlfd0YyQhwugf3Gr
NRw7vF8cX3ZtoRmeQScmsh7RnI92l7B9GWxMz8uWnfx25nUK2t0VBwy22v5iWtlsR+Epy0fV3M0r
Hxndfw/dQLEptxUSwd6JCNXl95082mC/eLGyHFhQ2MZvlonRfImUf5XZLPoLG8Fps432tvg13PM+
SMzi88jN1XntAETUL7znDm5+GoDr68LIWkGsx7D6mNnQFEn6aWgUZ8Up3xTKIeKSsarLKXzpYt8j
8dyzg6XdMZKy3MgbEJVh4Zwj5bmcCKxyYg0JWikARph1d7hi+B0hRB2830waqEto8ijlJLUDK4Ba
9Ju8rcdqiWknfLrV24J0UpyrSnLTq8gONaG/o9rs/XekaKIRtTYxExSt1Ek6s/Hc5huJzzV3Doxp
0/q5pEmUB3uu/iP7TKGKX22xIBqcvaQ0yrzZV2GbXO8KI7vJQf3gpALfFUZDLPc2jei4No1tbyNo
UDzSUrWgLi3pPz6OoVM6liu4ZEaQ0CiZo9rPrXkgqrKPYfEsof+jYKHLHxzLvozD44kSmkRwGQAn
weCW+0+jQ0vl9uO3DZ3WEQ7d8DeMLsGUNiP5ttbYOMBlGfjQPiabiJJZBIpq4lSsD0KgAP4SOPQ0
muCr0KyOtbAhhy8g4mKtvkta7kcql4eKJZH33nM/WVelpIicQcsNFSijjFKNvWC+Gvt6bZHmCK8k
Ifl5BRUSSmPEBiXlCVAc8y7dYBtBPc7029FMoEvbLkqOjqjbSzmyGY8jRd2k31J1QPVXUV2zkSXk
QJu57kNaDAzEWhxTVBYFUyEH3WAacS6K44Zg0H3lXYHqVRyY2t/XcGwZeWlsfm92k5SiFvzGL0n2
kq3EWxqdT/eYZhmcc8/sRR0D1Q9Ae16It9ZSvhQ8GBmS9GDc5keZ4c+OMABDm/tCBgyNeiALo5LB
+imWN/zg6Ae+iYjTF76ufxrOGLxtrWxqzM8QP45iqz4LARX43lv6dyMt1Rm3XEdUFsza9jv2ynbU
wzTUw/9NcBvR1jidoKuNCGFmjVqgesXANNQ7o4SapUd9tYyNt70KiiBaiBTfOHecpVJhTrisT+o8
uinNRpdMd4Y6YwUb218G4ykP7TCBOypgHrV7xPgA8gIDkdB9LuWnB8+/ePwYN6iuzO+ZiXbde+uF
f6Niyg8Gq0m1s4R9Gjuvb8dbe8N71gcxkq6eH6EOovnYPrjaPD+G4qgv+ljqwIIcxfjmLEtnSTeR
oOf4KY4QF11ii1g1JTumZS01Hrnlbo9yU4IyU0/5T0+UB8xCz7w2EaJdqV2MPRJhMeZFX+ofhy63
qK3skFHMPwy0lSvs5fbCTwCxlEuBLWQG4sz/gVzy7zKbelSQaRDS8w+z8eEqAfBz9yo5v+94zolj
zgQL8OkVltDEC4Vmn2SiHu1mZSF9E4gg7WkhXINlQIu34i8L1bYTyKEAYxqyyzgp5+OWSuGkUCos
FVQhjhCzTptFfsKocs3cU4c3jcQ9bhQ3kmNtdUdORmLwMiZMs+Ikei08p0UcIH2TCdXNn6weIPUk
VXduXsOO5Cbl1HT1EcKtcYYehD1hUvnPKtR/04XLoqaSFjhvRtXAudQ6REb8uri6IYf/rCKVYypS
7YWbtphvpmWhfmTxuxnRtSYWlMKKNBnQaJf73XABBszV50t7aMinkso834OgPognYfFHYGIDX87d
8FJK0WbYlFyiZ2e1PdZpkYR/ce3s3bNjvchRfybsEA7tya+5dkkmIRnYEwS8246Woq/0BtqKx3EK
+AJXOMroGgBiJqfeAeD9MjCOMjTxCi7HXh+2xMN46bluOdOBHkAiFq8bgF1M8lQJEf4oQ/YI9Khn
SY34B6aEef13W+l2qnNlkcs+9dz9l1qPuxKXC6fmaelk+AVQoazg4XmViMANAaI1Vl/ap46SrfoV
hRovO9zuWiIL2xNVG/G+WV9kcB8EkzFz0KLSMbtZctWc3FU4rErbWoKm/BQQcGGyN3Z1VgZtXXj2
seoHW0K7k4dniU1OTToTQMTIQDoru+eNuoOiQPkAoJaViI5VyWpQFuv17cCRK5JEJjNJCs/YwL3A
v0qB7rTbVcZlzr9sO/55rqWfLNHVA9/zArCIHcmp9GgZg4wJHrmrvnJ94zZEmH7wrd5Jo5w6F85D
7uEFnubKPqri3MiUnebik0bKOLUqYlNQEJTl5JZ2TrGPDr5uIrsAdn6rmwFOn53XRQu+T4+qCKCy
7s06ezwaNmmQcTKJvIqu/BwnVa4XZk/a6JjvN6IxAiMkf7HMQhg7H/KAcpjx9Lrn11taF5MLAkfl
Mx7F1X4gOrpSUpJcJO2fCUlS8EvDoJNJH5qU0X2taJ3t2V2jO4k9RGWNQUfFY2yQ/Z0HUiNI06Ma
nwd2MsvX/XoVIxsIWW5wpVgfaR6SedRd4d1OxXruU/Gg2xM7CXno7ma6//p4PYb/UJO7XvA3SIke
MHkF6lmnQ83jXmHhySw0hMLMC3hBaL0KpZlFp4uHAoGUPXacEU3ctRkL46Frhmtzj+wA9S5THMpr
uBhkoiMOC1tROpYbpr5ifqfJadr0jUWM6BxBHUQ5HNAj0pqEuTH04lXqM3dj5QHSKx7YE0CVVNzJ
6ifRDDqroNXpYRbQVmQZ2W1JfJ0nfxVEBgeKF2zCmG+mM6PJzAvbQ8J6lCA1vq2cRC5qMWXHv5bV
QU1/cegdQ2CyxtH1xQSzzYO074Z+A+i7D42MQo1Fu0kNwE6QTJbFUM3FRT8ErWim8pTz5mD3DO24
gpL4D0nW0jL4IpKALSdLvIeaFbTezmUHVR1mbpKIg7R6+fa48r4hSkeCOjs1nST+xpC/hfExFnU3
UsTXYWGmaLZBHg3XvV3GFSzabmHEoxCFrxqnTlpk4LCHTHfgy5u4asuD1qUY0cU1RjKW+cX9gzt0
Vy3/N06IxgvSYxhiV47UDzAgvYvwAyd6IGbUtY1BKNtFIEAg8cdRSaA2hQrvVfwuU/cTEDNmH6xC
iYGvmiYErkpQ29UWccoZ5vb+XSaV/dII82yLKzGzBm54uGQOHth0qUEfMb4ZV/i09Dx0Aqvw+WGF
K6YxZWHGgZMvOWpcCkFbiEKvbeKlEnxWUjG/awdS99uyL+FdQPfyz6jq4clmQ8zI8LNeU0ICg7pu
zNcUnXQEQP1Lr5TASZIfQqF7mSW7VQcrrq78Mo0k2K8Y98y6e4WE8MGvMjxqblHy/Cgv1AJ7jY7a
g2BeXFAwjdOOpIp5JBZJrAaB3zhc2BijC6pmJ0R26c4A4sysafhi3jxMLJHxY2kclI5qUrSTVDSH
oub37OBDWzSJpJLbehJ0yst1Eq8yctBNpJ3bqkdRnAYJ9v/8V+fwdGntboMzpP1rj5sfn4E7AheI
NK0tto/vDS4QwfPip2RQAONSuEoUonBQsr0FJfvknKhV/k+DsH2jQkb/mAce+YHPQZSx2xsBs5Iv
MVkPJSOa0x33FsQJEfBCa+5P7VcE80vND0F2xOh53g20OeB1MuyNZIZwUTG7ResQyi9Z5zxLn59E
MRFDy8Jn8Q1qOxDyo1CpkWELYge67aDf17Mzgm+hXHgWiZUgOoIkf1RNdjEBtIlCVHm3psTrFu15
GWTc0B7Cva3Pud3Eaw5mxqsjEf5EssToxG04FnvCRybqf+7HbkWhtSxTBgXwXgjWwr5YPTRFPPwE
nENGcWQ4vB7AgI1WhRK6lvy2d/DJC7dXiyMm99ecsiY2wRcXmgm3VxEFMnJzRY/iC0SOjwCbzCF9
4SNlQe4P8Y9pZuPA4Ug7FuCoz2B6J8F2+jCJoBS1jiv+4tePszzwJt0MMY2Z1inmgZFxTRp2i8nH
2S4g3mVCBW/4eJIvePWAHrKUy0T/xei+hmBly6gzVyXDiLUsYbUv1AkTQVy/7UKmVF7PwcjqKaZ0
vKCC6Mo+mveRXMNk5cxF59J9/OWQPX5Zb4Y7A/lAYySdS3Qd97sEVWb6qYxM/1VBndmpLRLHIVxi
kiboAC3fO4i67JIbyxKVE1acMqWRq7qQKgBlWRJkG7uEdPIOEq9QFb55wep/InsPq5zVBfngcoEg
KH8pg2guXs9B560aSdEnIJrgzgzanGl/jQVrISdo+ffMR2322/HIRAXZQr9iCIj8DjeG5Z2GmMbM
vAGoermer3zbzFEJmO8TyrVcfuf2T00aQUS6G37Hinnk2y1dFkASyh3xrdmNSGGdtKZl/vj4T0zm
LeJkiHvoGuGHVaMbXvATopKLUzvWFkOOj5IeKk9XO6++q9qxcX20lG/oW6uosRX1PryBAtnc/AW/
J4YNEB6ToZ+9X3alDUFwYh83aW1RpHNW7xpXXMUXjLZuM87o47I7+5fQBtwhJPm94xtbXbfT7F6S
UIez40lH3eoRybko+YzeDwEqgDBz13Km6mINjDXcLNzZjPFV0itWVbolIGmG8ftyWBzCB/k+jVbM
yuOFuwtugwJZvohX9dgQwJ+oV39qC51UI6kwjGEVzrGFShPt2rFNwsPaQOQ4PLbYJ4Ukhs/Bm95d
IfUG85K6EemddPbZ6o8JJ7st40zcOVhI/KsnflBcJrMIRqwAjisW9Sll7mPCxxKClpsx6IxzB35k
9WWtXNR/xJvO2PPo6uNoSjtzcyEg2euTrb2fOjY+oporB27rJo4/PkkV6PEDbS0OiM1ddqIEIgZH
A/f/VKbjJAXlrZqg8MmZ1Jf6RPpzHYYTl7/eU4BUHN2dI2S5EnmV9Cj7tRlO8ury+Yh4uLuLJzIM
ytNSpDXqG8WODFfyxO1blaxfDFi42Stmy/KKM/I/Qur7z4yBdTk4vC0umRo64OUKRCGXuMDsryhV
IRzMcXN35TdN9YsXrWS/ouhVnexpAZp3fNPW7zHtsWBTPcWfdhgFPNMnDNKEitIN9apbgE2UYXaa
lv/fgEHQZVfFRIQqx6DLWNa1ZDJuZ1VNQ1MY9E2MjdYSn0bPXxzNtMTss4rp9740tjHuoSgtjPnA
80saRwhXNGPuO1Swxq9/HY+Sx+TvFexZmhOtfbcdfkDkHm3vQkhHkWSbGEJridwIv6iNbZvwWCeG
cBQCKBR8zvNY31luBszfuT1w9s7587a0DVDzMv+Me5KHAlirrvrblRFp6qotmw1VNt89ZZMzKYhX
nnqtfjmVEkz+tlvgQfI2VQe4b8h5hwqauJ7Rx64xj9iWueWrB4g63IY/ShP3aRHM3s9HB2BD4Us1
EEstqTO+/FgT+P2UHfdJPa+btpKiZSPkChgJAEbMt475Exj3Y8wQ9GMOfKOxlhvzExQLoi5OSqdH
jOMiUKGkyXo8G7cJHk1bNKq5L1UtYs7hgCmNnkmYvedTlcIpT1iHvmJw6ZWBWMb7+2+/2PdhlULf
kMuqG1dbh81+G0hXvq9+6xAhXFXxnE4IPCFhT4bBi/Iybc6PuOD1AWXszUu5iIuamXLTdgDU+hs4
7+y8YhHyQ/cTMwspy8mFhxwtCnLp16zSf4o+5drY3cSn3ES2zjuuMXnMjWdVSQHZQrk9CxxTi/tF
e2LyvnSzg4Uuh36i18eCvNARTpsgV07AjAw1owH5h9VWwwfApHzmTa1Dqu2PMDyCsH7NnhTjuSDy
KfodiBDeXADYtKZNEaThPjvC05kbiScz2ZUK0zh3tTuazivMqtNA/iyJ/cEu4bs0uYgw7aoj8PPO
x4b8PipbC3Qg5SYwBrklnuuCvTWS3qkeXj7LkpSoGIoAiPfY6TwSHxF59XDCXbnlHn2xKd5h1ALG
sMq0a2cCUgZDbif6rzYP/c/fu8/BOwYXbPmIUywDkIkYu/PV5uJ9aw6ipnU4MGn9Pr+Bdw3Fz0LE
DO/x1WAT4uc9A0MmrQ5cAYtZwlKi43yhhbUkvvUdW0f0GJ6qXb7kYOJ2c/HZaub4qbnUuhX6xPEV
BOZESSwCcF/UzV2glURYBOPq9+0aGWXXUB0oZKk2BHu3jiPSCa6727UqxZGBDpQD6blpvK0UDu82
+fa6ndAI11FHHjcM4T0P9YETIJSa7f0ncWGtfXOHyqeel6cUhYl1wwMuIiXxjCutfKoLEnjocjwk
hYAIw9sDzgtoM13gWlfBwfJwDYp7Evp/MTXq+9LL2lhETrufdm5FpJDOml4P9YxONrepgQrCrshi
OMTIgI1qNNo1/OLpQCFWZRj/B1Xv6v6xSH3jUts2zm4dMFiwlhbQo/ejdWrNBlY/+WADQSMis7OY
wniyWuoi7Mld6YQugYzNeyCuyc8JtmMxVY7QZlC6vp/NVUPQU0ccLkFYSZ4MbX0u2Bdy0TiQpfaM
ACIA+VF43a8h9M0f1ciX7inZMAz+Bp2Muung/ScLBMEJAac1cwTGssesHlI/+rRAkkRw+SgfX8/q
3lOgisvLc4ptVbQbU6j2hEt+Y+zpwQcJpw9Trg8/NUc61IgFVl7KglvpTkmxJV4dc7tOA1hprHtq
mvEm5i3rri3NVcB/j9qB56O764QDRztcKUDkYyzJS+vHSyNE8Zfwcg3rTtQyAc1elC3m/3LrGyZ9
E9MUJkK964yimXBcLdzU6sBwBS8n8RYTOnRrE0MCBujbJkxlSIlaTHbMPsL14b1F8RJaqR4cfcx6
b+NS1fQs2K/1vWlfnFg7rtvAA+1tCBvdWtZmZ+gdzdpgziehCug+L3IK/dBv4uixfLR1sbszbaQI
36Mn9tmLyJbqoGIl8bGhIVngFxYjIvXYtDK2tY3QjU/lkvNx9AM/tl3huD9bBUFqYiofhRbsnlZi
o943xv19x5x323er245hyBav8RXM9Hl4VPh0p6WjrQdYTuMhsH+NlO8BbsU/FB2EuNZ82FHAp77z
Xg4jdj6W6O865a4yQOX2eUqVVSo4efvq+qgOrt/rLKe8nsCVQQaOTMMFlQhKqrNWD+6QtIV8vD+R
xDl/o5R16w0l/a6lDUOhTyh0V1Yj29tegFz0uReWZLSxmM/gMceREwQTjKOTqeQ8YeSiF/wEokqh
8MNm9/H9aZZGxrrJqQXhi0u4QLG/yyPvDXQjD2O9yl7OFLZ1bEgaoKCL83kW7G9Edz5NAmt9KpGv
z5CIs8SYxz70JlHALEwgMQFvUH7f/ESmJF5uOI6lAs2Shc/cCSQ0A+cXN9rjeW7rJHCSorIMQWfD
q6LWDt+NBCSdVdS5v4nKJjtqCAA9Ma+dMf/Alo+H8IB2OQP89gvpB3TCEUwiqLR7sPcBgA5k5ya2
y7MRN4sKJ3ktSQYQ36bogh2fnIoYEuUjBsOFqv3HDrCUcfuMxOUCXJPX32YIAek3wqLD0GEjj86s
OOewFaAkICqbAclqINe8iJMeLGSj7xGB1qDO+lVgh8cLE/29ujcUqLGaGarCH2bgPaIVAwT4aUKH
jbw1PZ8so9GhUopNG9lL8KovFOXAeVK5yiLvOHRmY554Ah3DczEncDbwU44cd/+DTaoPPq7sG4aI
RtaBF9lvbqfA3XDBrScckYTmARbuqnA34uAPL3649GYEdhaJ2m78wmS+uLBeF+GxorATmlWmJ+aM
DCTrYzH4m/xVS3dG1a55/eViGS6HeIr737p4OikKqioXGDTv7IvbTzunleqH6nIJcdvx4rbfiQyD
OldnkjJYu/gXvlNeZFYJ2aql45WuoqCOPvkYu83Lu0CgciD0bL7PsZbgxCueeWmhVsJxWPKsE2he
3UE3krJv5hRUFBDFzKpHEP2tAgM+xCYWfC5xLrIHu9kpY3W94/7gld8001Q0p+JkfqY/QR5n0dzR
4HrruD2yk82ZmHLkRKCXRdtPjWF2ZKsSNIUGBaREH2x/bwuaqyZ4a0HnDheRX/mF8An5MWpxva4Q
8U6sIG8GsilwO6HvWpSJ3GZ8MPCfAU9DlbIo1VqND0Bi+9nImkfMuNh0Liu2pHZPqA/j1O0l+aae
Q7/OBeMP1axvCNPX3Qzhh551grG5d+tpfhP2bHAcPfIV7d7tRQT2jlcSrcaSipzgyqPyiXS2DcDK
f8I+7RMGHtXoIqHCLw4KGfntZgVDsaZLzp18PVZRYQTIXP0gccCB9PhV8nz8IF1nWyHJKj76+F4k
1ha9CsNpQGEutv7kcM21GWu26fGi3AHjg79jQJpDJnLf4mOJAwZbLRvFW7lU23LDojEl99665QLS
g5kjDJO7o3jqqZg4OODbyKvqT8YQ9eYjEGM9PQ2fLclxkGrSQdUXa/QYjD86j3Y0N2XSvXWH0FY1
YwinNfoKfBKZ4Gc4eV771j61kbsbpjVY5RztICYUgsGJdC3bR6w8/BaB21RWCpjO79zJdho0v8Q4
gRysZ72vNi8m6ZdNLMRP9CRymgvKbL7xCPweWdDo+BDsRJUxXsBH2ZyCNxXgoDpx2Gld+Z9ig1lf
feDkUceUkwNm+2VwRpA95O6ynfC+5PsUQd7WSyRwAOzZNnkeb6Z338hnaGmAh9FbCabVI6uNqdBN
vFta/ANkoZmFlJ/4OVaIuGCPhxpm5RaCFZMKdpdOAg9g4dM6u+9DqJPLKkjYZVqGYAuxsq6PTnz4
wCqNUFV3SkBJOlf6X9UUXo5j5Jbts1zV8CSDD3utoPIJy5hTiYcNAk3kdNLSd/5oAkgIrcqHRGO+
5t2d/WBh7mLStawICBxb+QvD4SCvV1BWE7x9QnoiA2idV6/9AlIk0mdLG/j4H7aPF827ZnA1GHRO
LEqbAw6RyKoIUJx4JlYtIK7oyR2xZPtt6KZCuu0fTsFGliL4FT4IsAywg+0zHDZ/IjOYUP+gfEcK
phcFjEae/5JXpkYLB+xkamFISYJNdGWtz0zN4Jqp2c8GrdXkFOqzofkgFVD1UVv7Y6+nYZYmLShu
HaSWgm1s/CrzD321+fr9DgQ70nLa6K6spdRkttyyAhEmsxkNaWp4/GZ5Wyzg3UbSefg6kZioKIen
1HrMbmsICtEo8E0/EbtXazUZulZhHlWUzrZoQEwXuxhmEQYRs5B73Lybnbiu0Uf4lHSTbU+aVtoV
jadMDO/Io/7pDU8HwrnylNhblEJyH3/Gh+jgt6AceBVlCD5g3kDkJgqxJvwhCKOE+Pc14HcTPxMf
jwYsTlbyLEqShvqq2agGqZvvwfpFHonNVoGdBBzb+WzXxMC9paKlK+hMxpXCuooUeLSid+oGfLiU
Z5Rz8F8xGaEKUUH6rtTXUku31arJ6s4n/mmICmptgnV6bJyUyu6hnZvklhPvbjACm2cWN+aqkR+E
lSNY8vqIMhWwGZ+E2765KDd+QYt54HGIE/lupzwfQi6t+vBeUtwMEr+P5edaQSCq1pIQyzSAmQJM
U6fmAWX8QoxR44+ayhbqQlt8tQmq9LYxPH6wwtZp3M++djgUf2nN9WxoY85WF69Hvzr0l+GSMA5y
n78qb4KMkPyiBKptlblF1cA+ykEtyQ+UIRh2qr0tvZBouZRws6AhDuAKM3cBQzHz5tzVZCN0RFir
SFz+sitJhXV7hsiRXvEqsOT/wLTbnysw5QgJU0ngvhcEeZt1+maQKmJSObxZGaO1AxJQYCUkFEEj
XzkAUVmOE+qmeWqniLj8T8NEIjAjJglpqG0ZCVpu8ab1OW0tfK7jRFUz0k4g1vicBru6HMMJcijT
zyEZHB+RsmJtqnZv63ca9f1jncRQyqiVazvOa2wPQ5+3zMfwc6n0xCN7r8KKc+9RtIgi3QttPLno
4VOwtkkHXTIEzcz54wcxkBH+EsLoqt4Cc5eHPLEwxs20xw9e8Vu6Wf+bE3EUhIUWyLzJSGS5kFZC
6K7N3cVsZpTlQh0RpjS+R9hrbt8LiNqc3Cqxplue9zExmVGaIfhvqbaRswe/8F18XefIQ+b76cHF
juPV//C+f8Yy88JBMegcNPmQpdEEtgyneiq314PfeuLfmeHYe9HfepSwKpi4pwRmJQYKN7pc8lS7
YcFXuknEvJauGLeiULyTctXuFy7E5SPrfO+d/FHziEs3WUj+lAQ3wIQJ5hx49JuYE+B+Pace1v5M
UyAe5oh0WhSJnE5LUVImh04PGSpffW+A89DNb1xln5RQVGeeLFcKFOMbqN+rUdijwu7BWAP2R9EE
w2wl1dJpe+N+obhczhdaB6T/rILZhuLY2ggWDJGroZSxx+mFcNc8vnWIhnN2fe/dbffermsWYmK/
C6qTtBmtFDxXJcm6e6sKD3/neprTW471Bket/418VbAMpBhhlQ4LlhRcbVpSMlf+TlZkkOgw/t8r
syajr+8srU67MlBtN4K8xBsXOdJrYd2RCn5K1i0CFJYAxnHFg6iLOcOMk6JGBqLpMrrWfWK1TrjY
IoCIZN8Z+/FSzodBNzszzmm35Nmjq02V0h5RgrA9zIFFdCBRjQ30Frg9pP3G2co8rPWqx1lB48Gy
LZJm+ewrR6TN6wbq3DUWI1raE7+M6zZB5TB95s5Y1nAeXREvhOHYKxjMV++NIyaH4muvbUbYumom
7L1PN4oVD3SSTQeAOoMKjjN0KpldBcWDhAdTuBztDyURnWgpKy4NQcyg2eo0gbRgNQluVlRE4qKB
F0eCga60qFPwaAZ/h33mvepx00IJPHc4Di9YmmGDK2Mqc8FxSxdco7mu5RUcdhOUcCpTK5GZysG7
/lU0BmWWvez2VqNxD1LvOwkT80rYmfEz9JhDLktaOsdmlLHYL2maVojLlbCzP6Gcq2eIiKmyfK3Y
8V9oQjERSsac07VCjLE5PfBnrYRYf1jb63/qz3Nq/HOiOAP4ylOOXfviPsDY7fW/SVg2xvasBqw9
QDACbFb1Hqr9PVwACdIAHU1EeXDf3yw1M3nCTqEcDCgARRylBcehUvDpUQOK+6uYrg8a9azmLHi3
vRSeY5pk1hG+2PSvt562t23FvOLLbcxfcNEsp8rCBsnEmIQkaIopXuRlodU+dgAznC1xkhwOcKU2
QRpYSB0WEFjwo8MIOViUkHQEotOp5pOCQzWnjFl2sDD3/MXZRjIuMaKUVybuVYXSSXyF2Bo6mf/U
r6/ihqAeL6Gi7zIyRLMznKcwTABW08whcPLHpACtNTnxP/t3vTMFhL0UxxcscLNFghbkefMAXPMl
BgH1NKz23pxjlm46AZAF7G9OqKLl6yoedLorKGkOAEs4j1W3U6rK3RTYtm5cQtbReOTwMb3HjIRf
aYK+CKgWmn6xYQ5dbMFF9iyYgPlMDIU=
`pragma protect end_protected
