// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:04:23 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SSA4g/0wQyktNBX08i6gXrOhyFUN2EnvOABAXxZ/kQ5vZ27eKTCkcAzVtq2gCfau
UloYQkmYL5RGqTEEWRcgSWaoGkeh07VecBnDKHZ5ZK8HXJz9AwLEV/jmZf4hqfKP
13FrUvByedp05sFcbOI1poqA3V1g9Ywoe6OwKnqz5nQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1760)
DannTPoMmvGG2PoqRnJH9TWNOqymcWVR6PfuswgY1+gpagKXQbJWKfYINI/5oXZ8
A440gXI2YI/s885hf7vAIwdDs3/phRC4S1fA86uF4NRTQ//goEeiKMuiEwad9c1k
iL20EGgVGvWVg61bAT80NymA41cEL+7TSBSldXf4dxDsu5wzrYh2XdWLuF7F8AQI
yqSB8cxTR8SpktrSIthd/xGGeeLOa7lw7NN+6AbXBcPFuJUlEyvS/pYgtl1mqtDi
DfQAZTSFmTaFqkLbdMUDFo5bxwDS+uHUv3KZ6Eiwptcou7olcCfoq7oOmrY0+uvv
HiBmvtB4bJXufvFGha4ORZ9ZBLp1hUt4MrLDuG8XQWwPPD+dTWlcqRa+oSfPzNoF
/nocXjsTm6ucmsgDSiWzTGfuQiLxf3/kRM0i35DFIsDZmV0ttYOKWCpXO4yutpt1
TdvAnmlSl20A1qpppRyRkqnfs39zKplrCoAYqisxPvbVfmPGR1aa8j0cccLflbTw
CeCmq6TTc+E39HxcE6ucDZSlq78be2ulZt6sVb0xwP6oqj2KOw++2eoOOxGi3rXx
N7LqHHnAjKdjIhIbTcMtnbO21pZzUxQ6CWprng6M3tVHkGOviYjIoRiYHbQv3hpp
hxWqLcXNF4eybVANgzJVRDCfzfx8kfaOfkEZPs0hN1vR0Loy2BP8hNwyj9TCif6b
As/zz+1+4tls7cM6FJV1iuISgOGpvbTz5ZU4bCNnKE/6RPrdpBa4FZWjkZH2POds
UwdAbeaHU2qWgfVU4nZGMVJN71zOFe1H3f7MLLM7iJBHJxUzJdOj9bei1d5DZ1Y7
QXWgfRIH6Yeb3MaftGc7CXxYxparcFnF4a/jrDqkwzdrfGiM+XVmuhijvBzONMw+
istAyq43MetMVje9+OER6G75G25tX8b7n93nQNu8TqmIH/dqS7stO6WszCdVANeX
1tSYCW/yLbm3EcirgnYkMwrZSUNjSvxeUV2XYH9c6xJgvDEnBZ8I6vgFS9qJ42hF
1IZD6XtVB/4mhi+qiXEXQ4ehvTr7e8dV4h9hymSJwlbWOZpGMBlhpRhMqCUPZpqh
jMbKnSBKvZOeXIXdXffYViaJR7icpzybI4GxfH6Gku3qVFNqcoHRJA+h2UFaR8nJ
2H34AbJlE+LAqO3q75bfsrCN9+AXrLS/ZFNZ5rXygjTh1dZnmowCgYNctfH+K5mA
RdCDNo6lhe99mlhqGmnxAutp2UeEmajMnW3BgQQ55Vwc2UeTYRVApWedog3XRsPO
WF99FxcXVGyC9UX8Y9oFypF00XvBp1rG+D6ZeP97BbuNROPZsP5sWDed/zRIWXW0
lBPCP877iEiN8p+bOwGri0+CT4maIw0H/1fcLZbdDUsCr1+Rzqiwy7SyfvypYiSt
llOJuQYpjiiXnwlnW7fFuQ4ugexGBYBpwS4PY4xTwC2sBp9umrgl38MJljUAtK4W
X+4PIxa9sMDyyhJ7kqx+dRF1t3kxQV+37Faj1yBkfOBWO8PtUY+hQOorCpatV33M
dsHIQ/JT+2mb27nc6o5HErvSylvNh07PtefxrukFT7kQ8Hwck31PtOcPydsToX0F
x+0EBYytU29wnUxhf6eBt+pwEa+qV1kTLpYSPCFcNfX7nFj5uMKPIJj0NXBfis7l
61HIj/4py5+89YJGbBlBcaOV6w5EgL9ERvWcBu4MGjPoN0e0P0fJCCJEOLNlTULE
WAp+DtKgVtTWhEzgrLwIuokA2G11jOko3UMF8AM/C8BOTvzzKM0CXjOAZzXwBRDd
uJOirK0uRhBgo6FjF+bkyGNRT12BzAEoIxPZrzqOm0CGju7YRPJ8NGNQc/WcYij6
x9TVmWk4rf2Eza2IvGQ5gKILrYsJyefiy0dsGx9ksslJaj/AZku2+4Z3WUxLtCHV
9ChM8DGo0r7X8hU41OUg3lkHiKGK5ZFpOHArkyg0o6q18KlSlPWWsCtAUVR5RUA8
mD7EOu7uCp57s3K7lcBkJAGp2Y0uKfCsLCgNmP9xb01yN4HAIz3QOFiMPQ5dKmHF
wAx8cpPOfLpQcJ8ZQMPJjE6446HI6OWCQ/dA/m7A35aaNvo1t1G/duwU6t1Xc07Y
OUADNidaRyvznbN4y7EO6Mm/JQkwQtgXOCERQQVyy9hMhEPb4o2GQ+wM4csjWkKR
9NpJ/+VVl5Zv9+Bk2jlp3q3l8eTWUR7RTYlPozj7lAZG/wyzlV21boXu2x3ELFKW
ROc+7odBakE4eAvei7kJuICoIVZCI5jVSFMgKXav1rimVntN8TQs2++EDSlZ1R+S
nvFzzcvpXducuvXE+h2fCmMdKGk9Nzz8cIpJqx8yTIE=
`pragma protect end_protected
