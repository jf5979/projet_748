// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:04:25 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Hz88MIEV68HbP1S6BRZf0zJAYqPh0Szi+vBBobWea4/mYvFp5RMhtdOd47I5Hwn/
vCFOtGjlnwobVD8i77bhtKHFL4TNkM3gfiIL43XYiyXhgRNtom0TPL8IEIit1GKN
rQZE3UKcMse3DpT/S6Zjc76wZ6i0r4Si4FCXPJl6u1Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17456)
ukLBy1b6ZYpYXG8t5OMZ3lBZtxl8JiyjyU1WaCS9PpaWCimcrb+/1ksELWUL/AY6
LcfyF++6QEjL/6qcMb82oAAb+2fAm0i0zkGIdRk9hSDf3Bi5xh+rL+POeoey2+Xb
EWXBQuxpU+9rqSx8BMCp9f2pfR5Zh2ByoaE6KS5+yV/OLtmJVmmyqkU5uPrIzwQk
MLwXQwJm0sED+l3jW8ML47Wv01V4KYNuPQdyUVUTfx0b5zFylDbs4l1Gh+M7Q82k
Vko++yt/DT3wPWploPxXu6FZoIHNbFoZWfILNaD2GtvUSTduDSlt3qw7JB5P0oIb
1ov/F6ZWIVnuP6NpbKQu3JUbGd0osDKv+KYLK+IhbsIwZKS+bMxshG1jO5HiUMww
ofk3Rbj3Q6zK7w6v9RYv/Z+/Run/jMsXnC1+2IkKx+zk3pyksBje3+zQGmX2s6pn
yI+HhnWg9wzTp17dTg+3/sGjvHqjRa92BJYwodoCIru1QGln04Ivt4hlOp9ii9z+
DwCwUdpkR/9bW9lsNjP6WrsJZuTK90NAvuQep92C3R1ZnqQiWByXR/8wA0wlJXCP
D0IKcWNR8kAEcPmwsWdYrP4U5DG//cNpVzxwqgvk15KsbHY9jWwzOilPuYhcfEdr
gC0he9Emb1BXC2urSsvEKDY9BpalrNdctUj4A5Qj+crbLgwP0B3nwu24dhXtf9W+
QymMhmwai0aqq6787E9r8kKPtg7CsAXKr9c2QsGOpTyatQjN62QkAFn6U5RvJcfB
GmXWM+vMMh7WP6YoDQrFhDHG0tsNNrB/zgAJUJHRQfHAUFb+JJkBLDdfigZ/+cMa
28h3DKzNQpQekKGPUpSIyuIem48lbj3rYIKXcMiBmRdS4CSNR+lP5sDeC8vb8b6D
ehTW8XuimOQa607wMnvUGuDAp2oA55qT+R68T8QlQN/BzLQqawJw4nNdVIBlR1I/
vn0Bk/2BfmNuYu0z6+uD7Bgmu1POhk1DcU+rRZRJ6deGJ1xkwn+GZWr8J7nkpxku
7yaDyBz17xnrIeIbkVWePnW+jIbjnvQETW9LraHj2SIDvLVsv0QTmdKt74VLBSPo
rcYY4jkRMdz51Dy/Rt1w1J1TC6VmypA/UhokEW8b0dl63PhslExpWmbbs81rcGak
aDmv4AZ00NF2hNfs8+AkRhRocjEyZHOl/PSykg7Mrsw/a5yB1oKnEikVzZyEVq7K
vywQbk22l+fkPCeOWB1SBXNZ4686EFSV4lE41//XsKjyVsLBUXj9+D1Wu+B8f5Ri
c3ey5d/WvdI25FtXftrUhHom8hw1EtLLA6loWnY/F3ulYI3U4iA6bUBSfpGpC7OY
4UHoH0soVUdYNSPrUo7Ycl8sEalF1z5Ka/F741KCjLcWdW+GGbct2lKcskf5UwNf
YdbU95w49Q2S48AGfzIK3oD2a2K0/LwR+ZflMaQ8ljTMPK3TGEcvDryLV/7H03Yu
rx6BeCsXlaWSL+OyOfp+m+ew8ggrmj2TslnT0kb6P60sOKwkk7Hch4Gk0f72l4w6
kBqPxlqRruJ0XRDABx6JGQUz7AH12pqyeQIDYJhD4y6rvUbkQd4z6WnE82D4wAhe
KNOWfJQ+XSZpZRIw6iqxdC4oFr571YUwcxDlGF47Oh69DZXgiwVyj5a9GpgbXUhS
kvBe+7R3O0kYHJ5czGlWgAF5YWWUNBEdddPYUkDXZVqcXkVIAIBbUMs1P83PrAlw
/0ETVQ3WtZaBK0aEla9SgsnDH7ht5xozixQ9JSrcK+RPR56VIU0LrAIH0rq31rwW
h1IoVD1Gv5YWgZ+700LhBfDX6feL2pp4ieeeG7vwlo/JhOz3WqjBls6VAZ7uX9Pw
eWgatxWXxCzBA3vwCNR6pxOqhIZSQOnCiY3O+GLsqh5oaFXqsMgNrel+fp/YtexD
hVOVqFGH9eqh53Zhu5BSiLBgrVcAYsljY5stvBJiOFMmrER4sk2F8Jo+E2VHmTwP
iYAjZfLWbCAo48ddK1ZBFu2JkOLiwa3X4Wuwu3ifIJ2H5YHW5zum37Oo1M0gBtGy
qiNVgX5WHyTrPSjgXTF3kAi5anunql66urhPm59JMM4vs2Sb1kGERChvNwv5ET/X
Ek+cSTq9xNWimNqVTdksjoVhJQanzgFE9txWUMXUcDqDMub4QWK2nsJMG9eHzz3Y
zD/CN8UYkrDR/ZhCvaU86dwjmRDKmdcHKb87ChcMzqOaZf6JOoDUQG7f7Y73aMUD
WRj/G1n1qlmdEZ+WclSiXpVNihKsTjsYSTE0SkslWf8SrBIzoWoZweUR4eNDL7sF
XTSzmjjMwZ0qQ6Ay2e06y1Je5UlhEVPWXBHlFP98y3HIo7Uty2vboQIe5v2ehU/5
pHHcI+ipuSJR1tMPoQG8zdUMxj9nlV2noAE2hU14r21z87554Jpxe/iQ1QouYgTi
J9lteK0lP05F4IMY7Zg1jA8VoS1QEv8xuT1Q065EfeWs+mxYQz6fAaz6xWB6c5hQ
2k56sK9Aql5g3a1LLcjNiwE/sr0AlkqnUNJoMg/5B4qFj/K0SiI9XGnwfIKIRisN
mFxs9UVhPOaGRSQfNzQF+LoZujL+pz3+rez2WtD3P4gc82yvg8B1EO+EqGGJTD2o
plcBZ77ZklWD27wV2euGsKdJFpoXRY6BCoFstNVSen1yb4g70lpv0x1+IyW3e7TF
LBB738QaFpdGE7w9HZqS4dm+qd8qqG2TGRPVmTeGC9gF4HkWcKHbNjqW+BXIYlHk
yUsJvhsZ1evX62gsGd2jXbH2B6VtT9CQcHgp5FPPSnpdRT+ulBtEo3sCiLtEvZ1h
JzHs4fERoSMxX2zcGItNUv6RG4eKKA/bPtmorRxdvDIZNkLCNyJk/kiGZXh8HbUs
nkyZXIxYdE7C/JfocWbdKkP20kWvcPrRffQfdSDLLEtUD9e/escQOZP5gEJvjiPG
r9vEJ83c1JqS8vn2torezlFb5RPPP91NP2193MK/bvYeF24y51Xlba/NZL6e4AcM
NY/FIR3cSy+sFt387/1/5E+qnPoNPLze1M3jBjmto1ytzzwnYio5kluSaLDXyKrB
7hytH3s47s/quqGoLICJ/nFSX/107qvWWWkTZmFbr2WQHTh/n5kQ9+c7EUWigbgp
/ahBN3VTy38cbZy1+KIKudr+PWNJ4Ww8TJFtAtUEs74shCV3R1l5UiJ1JG0vQo2V
x5pe5VfJDdJiMwF6vandU9Hgm3qtekTOMIWWtuvEFAdLAlGb0f9OUG/P0boEDvi7
Pic/bLimid/K+qBWTf7Vw1zJPFvM92Eiu//mLcLQ5/p228e78iiObzJibxvSRacS
7NZAf7rHAJPAv5BZqLayf8oodxbLfCLS3eVm3qoOOm1gHSaXSh5zMtQlIrooRXt5
RonzNiaRcCbZbhorAceaJFvU9ns/MZuzZwFexaqQkoNKZusYWjx6jFSr4K8FE3Wh
84/Y6Ew48o3UAb2NohZ5XHy5s19i7WSk8JLkahhWEl1BOF19Vd9el6UA7VQzObN2
jxJfiR5noYpH+Z/8p1r3WJM5wy7GlJFHsUb5pXXNIElnzIMAeFZ2he1VFt8HR5qN
sFe7B+9HyR3BoQYG+KeFSq2QbFMo/ikCopzw6NhJbmmuvarDK9S6NygquudtrG0Y
JxweeNen9tbUgk/n2ETQLGzGrrQh/3BW2Cl9+ArhS792S42sZbXSVc+Az9tj3dy/
5URDMqS2bkgXZUXo2ynxGDHk2VCn4PH1JkCR3MADAF0UjSoOMz9tOf++vRIPEUzH
2rU+r10TCh7jpqe2b9mHIlHE7Q0v5lcpQpZAd0NnYjojiTXREa7SFl7x2wBOCTrP
N0odNbhsxH5V1U0PAaF98Kk80kya+PatTYUX7vvye8oSyYPWRyEXfBtvt7HHp2Ca
2t7OUExCayaGXkL/z2ZGCwfCKV0LmSgTi5kQpDiZOZE4FC2Xl0Q88HjCqsjlV7tW
YYTLZG2NkuDQW1pCdHDZZoUicbXzNK+6aoGpGu+kYmzrDP7c+Rko27x/tPIjmxV+
CGTkv9rcYJ5wn+L+fNDzOCDkMra0x+9PfJzIQnMa5A74l1uuFAiwF87vH8eo8enZ
nTEa3tsMHZfY+FSasVcjfDoM5kdSDS1IJhNSDhPrhy2FDOiT/zY7TNxs1ATUjveG
REkzGr5Cgd/t9E7RIcC7KFFhvh04D2OTYOHkDGeQQwC7ADN0y9oCgdrpLcfwBTqX
P+pYNh0H+CiGOPmGimh1hs8TyJUD+nBfP7D0hMqGWd/rlh08KMY7PZ9ina1Sbpkp
Dxyhg4HvNjN6qc0G2vpYkkS36i7UD3g9qSnxnDx+Aaspd/JymOgqNiTBmvsuaQ9J
TF7HJzGp+3JBPTx83nv/hvjRTyuA1T77UZmhFAqPGyXwnvjWltZS6E1AJNz6cbqr
XEESMQR50o4Rd4muXZmUeKp/M+l+lWTp5U4tJOfZE8nGDHrZZs8Hy9oWTO4XGvub
Sop05vS6UU1EeiCDFlBE5hk7xDeoOoetyuWJZETlD4l4f+R+JEQtEwU3z7IO+mRA
ttCQlVX0SDaFJPZzjV3TD4EvHt+9J3ONlBygZzz9LfCxKXXI9gVw7cAlvXDu/oPW
1U/lm6rH1L1If9XzEjnWI61wWZqGTGC8LLYmWQ6f47J8qiQK0M2FNInVydPe2ChS
brl3ZDzleHdxv6zoVFNjoKnX8LJAt2FoqLcuMbwqPmkSNSO6G67ifyhWakazm3hi
8wx/hBQ/aeH6VC7yxzDCE7itjGI/ZN03e68eah6lXtsn49DoQske432ZIrFWgLEW
A8QEs3yrZBX0R+ow7FBakliNIk+SlrL6R/fPnD3ITgKozr/zohTincdkB//6QUUN
PeeKR7Lm/iBKE37Jk03MHBafM6zl2HWDFdT5Syl6dnhgOilp1s+2eav5f9KD9G0M
kw3EsmPCE/BPADiOjPxbehszbCdpzAz6m4ovuzAN8BOesWfQrmrKmNqndR88kwhG
PHW+LBvuv9xFr57DmvXJqK/NDQlAtizgiKPVzLoJJOsJjpNgJrnQTDMxF/XgEtqj
8XPfSITe7fbe5q4cD7Cb+2VDc1swHDuzuQBIEhz41a15suKRg/9iZoqXROshfC9J
xftOiCQGCz3ClLgVL4wbUm32eiJTbgr10UIRTsVDSMW+mGNVVwIjKPGpnlIS8w97
lNj0jaMxUSFA6mLDhBsG4aYjWjYICb3oj4yxYF26YTQOp/yNXP65GkIDF31o8i1R
3d26pXdYckNEKGpP6RqVhrIUFJs1zrgRJIdT0kbl+aL4F9MFlHOLuTEkmDkqCq93
9DWuFfsdv43PcKPVQj9w3DxTDXNTBGazbfAfnN4fUrFVBK5/3eh0F6wiy25ey/V4
pWbsbP0n4jOyKzdl7k0/prpfPboXgcH/Hyn67nKz+HPaqXgeActDb3e645/7333G
/XLtjyfmndIDjZkt4VY7wMebwJi3hPI01OhXek83ikGEXbSL2BFdYl5f6INL+1uG
11HSAPNA+NluyEALVNNgOG1G6wBgGSrGaa3hXegBhn8dpjSBBKUepctBjMvPxjci
o5+BO0Q0Px/PR8x5VtcZzA0YOIY4Tg/bRdYQV2j0OVBTjY7OLVWAEAzu7Ufa9lCK
uueVJrqHkDMfqnCuDNGspL3qGNkr4pJO5iTg+RxCuzQjCii4a2iagHxQ8gGPnYxF
UCpXqMrvIbiuTlzwkQWF727kZZ/gJgonJC0QMhqUNFkV9fizUDD252uHbCMY15OS
SZJ0yfYcxEfza2iWftQ3hFPU+1NhW8ilQogYbH+E6Fy+4FwKZfTvi9TbqXpx4bga
0vc2/KhtyyzDqEzvJbe73xKxU2aNues2aZ+ipVLkVL5mocM8B/yqNTjfBPhI/KGs
S5q9AAXPZtpuwsgDUwN6jU0bjajhSmzRzN5QH0rUBQM2oYz1YS2vHRf727l3ckCR
5ZpifAyWLc9TyB9Cb4YQTX5Oz7pcSiJg9zXA+ueTYb6ztoWeQr8THmN8kIjJldkr
ZFd2UgIB3nnGFXvNsFAXHYOty0XxCck52NHKKXoqf0IvELV0axEJOsEl5eBR4AyP
ysBbw1ChhaT/NA98rNED9IK+ra6hsZzSamKqDhEtx3tRf46O4p+ueNvksoK+YCcx
QqdvUi9l0hp84YtfSxHzMEkYQ8x1trKCEWkQmpFMw/SZX4SfpdOhAxtCiEPBXcRh
gPdt9jnkYpUBFsuROifFokCPjNlboSof0jt/d0HwVMIWAeL7sXNz4JfIb+LpPZbE
wldT9ucPPGA8bOwh5jE10TN8JAECFuHQUldSTSG8vsNyXKXEGhN+n85piAGtdoFc
lknTCu1ghgCFP1TSjnBSoBrnhN4kB5fDcJI4jL6PzWOx9HHNQqGwQVNb7mubaSRM
/afDYE6rhRIiTUwbqn2dT7fudFUyykUN0d6NbkHRd5m1UThJHGSVudyuHpuiAaP9
ssmhBTqvYewrdXwvfbYtRq0FnSvJKqipEzX5dchFUg7rti61Y3MrY8BIrSktT0Au
v/mftGwXk0cxLtFMkLngaETRcykUfE/OKhN8lo6eRE8YYOnC9ZqFBVk4eLFxYU+A
mlEWFkAJoAXv19+c8nwKGpzXqYJZ5uErIrUsxCK6I4/YgeYuNBjQnZAeVlkqvdXM
wB9QN1xXuHkqQQsQUlj9ZcMmwcWjA7D3/yn3FVqT5c0iXqbLqpa2JePliYDpnk8T
I+Oaez0djRtCBIXy7AOvPUpCG6BAAuxg6xlQaL45l6vlDFXCmaD4z/odyEE3iIR1
NQO6P+/gI2v94FycdNX+MX2kfXv3a4rtXOk2Qqhi8vYOy5IUWFadkHZbuii6SeD4
E9rWrekqYDdXgDq7q+BtuwhPeWzolUoLzEvIgs1uTo/jed5LR7DFkBBijTlBOa1r
KKwc7Iyc86+yQgDI+7bzBSh+WLsefXUCiZBBwwwr+YnVW1J8l+LJK4nTmn8m7tUX
ilJmQkDivmZ5ipMhogY+bQjnBU6q7Dfm0vOTukY46lc7Rf2KzqbU3P/aA70J3Cfg
4tAXHFe93DPauyeceTbbeBiDM31sdbEqZGc0RWD+oGB9YE8BAVomC/4eZ6yaMd5O
RSuY7ZWOo2y1QWM57Oz4vP56o95hsfwZVCdu2dDyMxc5ltyqJ25QBSrqE0hPytLR
HxJGA8GBitpHgjlsG1oLh86A2rCKahyq7jxxGzIzcolTDb+mbiR6LAUaEzmPrRPc
JnvykDKxsmGBB6d3TjUEH57ocb0vBJydrQ4IBSJO5snxMflQetadiAoTAtCm/72b
yYGDMU9HXnXNYtiLe7EmyxCygL7r9SwsKm+Bb46T86TLD1fTwYkgDZhhHJeS2wXt
vJ4GAsn5KFrUs6511j9wNKKOEa6Ftw9tfrUmlbjz21HeD7z7cjyCat9MqlzeO38J
i/Qa/mfIHpnQiqvxC7t0Olll6ETNvVZqH2wDY5ffclqHV/qdMVHZcu2g5XpWgJ3M
ZEDu7F3LbtwxyXIvET4FIShF6Je+TJWWChmQArG2qP+8ehM9ym5sAkgBKJ50xWYT
z5XHqIwC57cfV4yzZb+/+BcSKN/tzRZoffAZGEo2ZI1nk2mMeALGGp1ZMzRqu/+6
iki3TRBzW9I7ZG46rdh+OYP4m+q1NblgnLv58zvzKPM/EqOXaGU5TAygx6IMoQmT
oycCTJN3tZhVVXaDJSije90uthuIpe+0o8WbjICyCPf4kyvVXNEUmYNh9VtcHG/m
3UYCPIR5gXv4RMHrTqzTT7u04P/4gZGT3XTeVLiC8vla/5JuqP0Ue/TaDHP+Gmuo
WkD7fmHKYCHoiRBjwPmSrWbYaXinbrYigatq9CdhprecpaXudRW8bgorDwJ0VdDx
/TeDaw24VBWlELCdKLn9cdIB9B2SNJnTcxkypKH09LNb9R/4pciijB0AdJfY+gjQ
nFLpVIkGIEH+kDF5p8fQdjS6xmRh2FMAy/+CArkjZejEb++5PgzbV+plczJXgU3c
vvGu2pHnrw7qLRH2Px+Pbl7gb4VCU9zAm2lfIa7Uy5OZSXyWGxm9o1gAq9uijT/T
utyb661PrTHfAXnDHnDUyTuOefHzbmTN19wFmCLn+LSWFlZ2ZyPSMfosrlBnklQx
lt7k/Q0E8ayXLjkOGy+PnFpFsMmIdvyopXXm3+sfm5YthfpIP6lfZqiDrCmc8yI+
zXMGpvf66ASEclrFr3fguqKl2rlYjmFgtRKGP75IVdkI4O49G2clfqOy57NTmxp2
43cTMUxhg7fLCBE21u4QgJ+jrrJv9JjvY/RFNMK08lukZx36PSedZ1VHdPZ9rUkw
0wr5DPDiemExzZN9zPuOstwQhd2OtdN6oyKj+fLV8cVRQZh2j2AoFkG6iwo7CaGI
aq89Q+H4H5qsfE+fxY5Ei3P5X5xf6gHLMRR6wdVo8koldJE0iKZGkwY1EZpgEot+
eIWrRDKDHQ8kDIyiRbT2w6EiQfsxJKnFVSBctslEOhm+XF6RfaMhYRWnSDp3/qna
x62WKgCuBpwFM0EK1bU4hFW5J1bbBHhVddKOK7FlVd3oWi4U3Hd+vNFo18dX3gsv
TGH4rQp9hxzfaPuVgdI+/n2V7jbx8Yp/YiZtbYafrqqed9KTqanG0NTCnUGjGBn3
2tEIxjEWzlHkASwZLJKgv+emsco1ZDs4rVm4Twrwn4EvtcFuKmFQmrwjMG2gVDrb
Wd2sG9+O/0YivKksMySWx9sQMyiKB6woGLnnfObWmaDk3FA+Yeb2BoR5VSqGJT/c
OeaMc7LQXiWmBEl6aaa9GXOFPX74MZPw1gcaxpg8lmpB8S9jY8inFn/YeDRZ7CxH
7+4P6h53ysHJ5UFQ1QUrPbiDiwR45xxMKjnc1vfXgQKmwjQa+EEEW/IZdDQ35wyh
0SXpgbjvRVBnU+IHJ0MV29FM0rqDJVnM5wsKi7xuzdXCoyOrB27V8jvBrS5Ikp9j
rJWwPP7rqN9eA3Tew9qVxl+wwRy1J01YsR4gq7pKKtVQqqXZdFsW+gm23OpZC2zu
SnHFb4C01sMPs9Gk5qXCTlv3yPs5bYJR3r4FDYi6pMjIryq+1os8u0xWriwcHMCn
LsqEDadHxJX08Xh6BmkuY1AcOy+0GEK2rqnDf6K0sYLYNmUbl79HhTdpb4elF0JO
gl55t1F+LxlWIG6jLpBvo66ZUlK8oyT0ZBArfigAI7kyNTzstTLnrtuuwuKA80BL
IjqA1V2MSD3PbUk/00adgFJNvNWzIx2yCp7CG9Stp3jTKZbho5PGFiFBy01mEVYx
8tXUqs53/AkpV+djuDFmzlOocTsQVzLICd4vcgVOIgXSh96pkCcSY6nF3GoO1alD
b3u6pXY3gcBrA5WMaHHejcL5lgDPNNn8sJDHgPaFplbTLs8gIPQZf9Hzh8uEfU3L
hxPaw/+CAH0DkabcbOjMOwbL0drDut0JZWipNJyCUM9wSgBHja4tY0/0xZG7VR7+
yju3hU+aeq6L+wv8Pn8UM2ylUA+HPNwLcePLTP0wZ9N9OjC7kmwY1BzGUBXcYCG0
7FmeJI0aIby9RopGEcF3oQ7CxW5xGSvsUIU7bpNKr/dgQdPT7N1YTmjeEb2/P9sY
4we28vH+XEGsTOMKZ8nOZDWllj720KthHjgkoR9GQHZCVb+bc5bMTtC5L5zVTOvH
WXqe7OAzytnSEJvVGrLEe+SEgKdvGTmXswTFfldRh6LKvuonuSJ2uZ9PDFe8G6dW
KaabtUfaD3gv0eOkuQqBX1XGh4+Rh16sbPW9DMeW8llsvK8ZVLuMt304Vw1mXOOu
pzO5OEzpYfhhIK7Q1aepg6UndhNomDHY5Kv3nz+5oEM86+ygUo345x9avgVte3Vc
efgKF8NXRUqDetZQc/9SE8xd6e0ZVptRvHnB25mF1JkJnpCDHcfdbROL4S4SZRiw
xeOUVUqDVUcvlyURV9ukrhq8S28d6bA+XLxsrwM06Ty+43Sged2SVDjElxkQdjmF
fPD7g1ffsjEB9XNzkl678NZStwvPyYtTgbiQVNXtQgnu9xnr9KCjNzFdU1yAJzFw
PSCb9OXzzHN2/2+h9owLXK7KvVKEViLqQyZiUD7PAvkkieYl024uhwF1X77Ra8nZ
cdeaSoRr3OZzCvMyeB6V9YelDz7zVAtvHEU0nyfNGZJFEzHaiv1EhGQBKep8Y0RU
1P39RJRiY15H8sdbSXBVzSjg8sxh23QnOauOnOk5m1KsuYMi11c1Fekz1FuYTh9b
glGB2OFqwBDDgXXc52QzwaYDB629UXF7CiKGV5hqGPThabQeHAYMqJ1kRcp7iibO
C6FX1ZdoXYNz/L3HB7dmTW/1SO6IcVtgUL4KqZPiEepPjoM4dxUwRXwlNlt6y2/u
UU/w98hUp8QVHqFcQCaeh946/U1FBuv081EFuNLFMOIQRovZNz78VZq3vQ1W7Kzd
j0AVrfTHmO1EOFRDcyS8eJzmQpitUMAs487jmBiLMLjQYR90ZWkvgDP5koFZk8iA
CiEK6ruBXrSzvD5CMY+BjOGVmRf1PvFZBuPp3kOwoXOTEiFcFvQ196xdtciyXEQy
3TEiJvMLB//bZWjlUGomAzMI3XurgZkPHxwGKFz4iqMe+u1Ig3hrBcNNhF7pAaHf
tV479WELitlhbZ+/oCet5vswPQSRii9uVvigZehurCaVKMwz5uDyNBCQokpVtFSO
rhTclTBhrLhSmLTSpfCze2cb4yKoYK8MIYJ0ve8txGRdQSNlOtHSnuWxg9EoU0Cm
iAMjHHpvtJKYpq67R4SJh5xMmkthtkxjZfB4sLDr+hwK7kqD16NeqfI39IA0bR7g
+bWJwVAWsAkmQyiCcHkaKhKN783XJDX5SmjW05A/Y+le6fmknrw9fqZQO1wW4zAJ
ARwDOeTFj3dIYSSSTJqWxHCv0yJ1hgWw5qVWvbKu26cyNcXj84y8uDBNaQZ1j52L
nnz2GFbkSLaJkZhIKrbhru03UpMG8gJnO3fX4UWd0NH9uGekiBBaJ9gPng0Afrj/
dmX3PGZpMjQmIgicZzn3xqBdkPkaRZAmgRuPxcrkjeHzHEWpFzlpWlTAj1/bu9gi
p3ZQxuDuK0VBb/PUrEV7bATlvBnIKRsSr6SnwVs/asTizjrEoYAKtVUUffRXtA7Y
0yZP12U91a3TYSlAje4SV45DmJLcg6F5mteY5jclx2hF+OCB01JEhP1fP7PzNIH/
peD4Ofa2j7F1CHeOYlCW4GCdN46+2FrXoxio9O1YOL7c09Cg0ku5xHWXDr5Mk/uG
N03DdjQcXKkVlCfrTmTCpz0vAdC7Rdd6ZotRmflwSKHhrlip+pwFtubd0r2qgX2v
dGsnLwV4vit++Th+ue9AKlvzs1XdY0LGWveOr51BjmuluYWelyw6idK5F41CTmcS
3qJHEvk/hu4MhW73qRZXnHS5JM6eBeKHoobMtVK4DxsvXM0BHx7d6F27aqGMMr5O
qj11Vr7eISXYapdC/i0tnyre2sA8FryBwLbPDMlNRhxQyb3+G5E86rsHg5vewNc4
XbpbNQ/Np8ZuIrVV0Z+whVyZEC3AyBeqMHWGGD9Pjdh0nIp2Knwn3Kr1OlTRgRe0
of6XPW5KAOncp/SypfTMEyzcQNURBZsHrj1EfgbhLrWixL5/a6ob1+TMHWbHktYB
NMX3b3Lf2KNdTMlbTgs5w5moDcWpMigzJ1jlWsf9i7CFRlXq1OpiV9n6ntJ1kUWd
2LJ/nuqeKXUn0+b7BJE+qK80FLBgqRcEuJRnViy1VF8yh8qmqbnu00E5z2bZwkhF
cpOjQKYu4OipWzara01eNrga1o3nUiIkr4rqbFhW5AlG7vEpSxYduckIVClQIhQO
B/2JCywoOwYZekekFFkYhk/+5gSQ4DRW1gUJqahQ3TlS94DTmKVE+SO5vzxnfZyc
6tjBPyE3RmTbKFytcmzwvaT1zN1fd3+UGOzVJrImBlzQ2XZ1c533lRE+faJPOoIE
a7hxVhGsw8aAt4Skf/jJz8cl4i7LYqBDh37oNwvRUah5sZv7arXMBKk0t8jF5gRV
WKbrWrHr3kfBmq6GwnNPONzVUcYPBWTXyk1yD6gdUtxRqU6XBHdr44Ikr+J9Bpbx
X1eSaa+58VGR5P4KKBf6UMbdcyZGIgP0hn3O+CjTg6fTPjgkHPk/J2s4nIIH5l5u
RoXoREf9lrVNCiwT5Fce3Wz5/dSwk1m0llqhBFTOW/I0jXeoI2GfRLnXi2BYmiK8
3ipsqerBhbfzFI+k4bq9tV2Z4VM8fbZYHTM6m5qsxyXQigb1QPa0yZG9xzJx4QEN
PSwrElpomXiDYrxNU+bxVRSElIKin7bTz5hgB59TpAQFQ07y2XpAG5Dt9POSyOlu
dVgTsS1myGjQwEfwfxjmowfrnWeX2F+hmnoV2s5qOE2dzbRCTicoZCrKrK26UXcu
NkguNuIhr2LA+O1kbfeFvw5tB9HVs/Wxcf1Y94Z/gGlyq0O23ZwBptc575iQ+mpk
NIFESaPLEytUE1U0FAspPzMm0OP/B5TGLtfaxNVLloCLiPwU2bu1Gah+V71lao9L
ftO++3fBZr9t1v9bbJ0ie9Mm0JNxqABSA+IMtuFYzrTNNSG7l6hLO1/KUlDsCfiS
ub3TdUJlMvB5wFGNnk3YuEe/qZ4Ds9txttyIN01QGeVS9UZUO07xjzc2W5b2qwim
XiKlbx3sfQrBPgkcxi0ffSAVDBzVYjJIrQHprljmyWIvNKe6fRYYFISz0G6KGTSB
h/TpumW3Aozdaz2R0YkvWvBam2i5Kv3kR141deiivx/v0NhjwCoqNKgGEmN6wS/p
oiI1LuUn8yzN9EDy9l5/LWaETwhAHtaqW2A1maBafWJdCRbtMlQRF22zDD9fZ0fG
JBSEn/aS16AKcNIGUOlFfQlYDRmr66zFbvI53YDR0jPyN5Fv+MevfzGygcvRxBE5
dKFfC/32dSDvJpDO+XZqAgELUMEpoX6W1TSU24gL47SRfbsariv+Ew00FtZhll7D
5W5EPXEx18/pmiHGY1eHpFEkbxv9lNZmfSHS3iCWF41aSmW1Pce4K46/kiPv78Tu
H+6qrTbCkVYoBDZuFZbcAspvHcvQ+4xHmPSTZ5jV7vLXPWomYvRCNHgvThRrhU3L
XfIns9vm9ge+G6VKSIvO6Vkdxv6qwnHQBRkn4BF4vYbzg0ixVwb5HHuX9ANgu/S5
4pAmy5VFrM3MJw87DgXJxBoW2mt5oGKhcjOmtcpI3NU+YN8EnnjtSN/Blb2uSjnw
Ll6dA4LMHJKQMpgML+LrWxrEjmY4vkzYT/eb0cXU3A5JLb77mgCdjZMn25GZwydh
pHqktkS5SMLK8XupF5PgF7Tt3xLIbqu2aEqW3sxeWq80X6L7lpdmZenhA9BlFy4o
OcNNVedMiYkjFxKQrsmEq7wEMcW+Lh2VV78jv9kGNg5QFrDgqJPD/FCwbkPWIDSb
ScyCasCRC3VmcVTiER+rLQ3xIyCsjRIy6i1FvARpk088YGwvllIorZqhvg7UsPxD
8y0ku4dxvGqzpOP7vCzXQ1u6dHTWwEvnM1/Q/m7US7blrgLDKlbhT7515Ly8FDGe
7kPOlZEXHFTZjK5TNVLwePNTAKQwR4PPG9gjjc6k99oOVf+q74J+IadIepTq+xBV
rjS3TySiBRDlpn0SUhKHOzuzEUOuCg/QQia9rh1cheNYKdgDbzwL8T5H2tqga2kL
QMczgI15LFr2jSHKNgFBT011eRz9fX8Udc6PQkZjpIfvmfli8qNshJFBuYIfdWS5
OW2EtLjQuuV2Y6SY0RAHPo82/GsvBh0Qym5lm2p6ub0uCz8/AZDKytYIlUA9mrnz
5WxLatNZp05/0lL5cZr8gJAgo02WD73BVHCWe/TLM+lxm/J0KLfWBHzXspX/hKul
HMqMgLqOnrbwjSf0mTOi4cPHUj1qpHDkNPXyGyRoWqaRfr3h2RJteeBlksgD97vD
5ea6rNPurJ55lztR2/IxfgcuZ36ae8p9Ry45Y+viaCK4P+lt9CODVeWiMMtMVOEe
87NEDFYORxQih7WTiD5ShEk719TiZD4tKvTuyv1XpB9EAq72geYUnbwKczBTP8ZT
zB0papJhjA3flrH0j2vgwCEPOVl3HTZJxVna31BSyk/J0WNhrBQD+MZvizO97Uek
vStLHXiHAL5fcAyxJ75MwfE+85LoATLYdFwcl5WiEk2zFKxwiAAKd0o6tQoYsBhy
EysCrDtLMiOHjMTuHIM7uTNP0yw984qqHf7rVG5oh1gbRIUkM5o+qBtUV7IAnV1Q
KFzuc0JUmh9zt9xxH8rsuTFt8fKUr3eWkPZgLCJ7++/INgtHE86LiIKC2ACzceJH
e6o8XIqpce7zfEA4Pm9ymrjFWT3GxOaDEyvivgtPnP4AL443cla7B0/Hg8aASNGd
0V8Ttdui5nh+7cXPFsc17c3U5TeGeds896ukUm3UVla10/kp+bF+p7f0zOjzh/SS
U4oC2R61nu9nYJ1STnz2TrGZsfLb7Oh3eaehfkx0JQWInFHv4cAsIpa9M3zatA99
QJey85PudvG9MLZqEi2noG2lPUJbu4yYbiSohPjQhB5wMTO0A1FZWDYzyDKROrwB
Nd0+jScgtCoVM7wedBZejB8qaK6CFDfXnTd5gvOMQAviQI877mPIB7Bxlvp3ChhY
vyUH8bX1p3s4STMDoUGQ3UizDdLFtaCPWrka5TLtweXcqF4e6AIFqbwpKqM8/Uq5
X3DPo6lisWpxwc1pOyWv4s59taffyy8FrVKZOxJ6EeRaiYwJddAD4tEX+JMcMhzY
Sj13MeYjRBT2EmcU+9rLGTbUY44ysxqDvHcO/Sjsxwt8UChECYoJLWI6pRUhBSDg
nrvuNQLiwuuMCDayH4uJF0wj26fjh18y0TG/Y9CKvCBUV1V2RdHDMeY8YGkWaWnj
Bob2G8BqicxTidrJnvfEQN49kjp2pXus4FpuJdANKPNA1bxNKJ6xzB6+fVvtQfW4
S7iULRWzijRosey7ND55XSuh6XbWfOnmVCRE847vENoREgByKs7YMYuVetXH4iik
I5LsfB91rwgmY6sb6GpoFPeaQGZ2skOzlytNxZuG6KCELdcMZJWyXxoJXBBvBXRw
7GN89azNfQo4p24/bfAbB8tTXZj5MUtoB37XPMD15D/7ob+0Wd4TL6agACulaXOj
T1BLAvHP5c+0ZmwjcuxTaAbtI9yxxHAolQZN4upd3y0do4Am4KIJqcxRIaGSiAhj
i0Cxjpf3avBzhPeCT9BADBadFzqChvquLePsYDJmnzRQzy4aVkeSgJ8m875Lsj/Y
HKAA5qTll6BSQh5sjdzWgrw23xuGhJptdRp3Of1mBUjw/jprZxTPzayzUdMPD7OZ
6aL3uDlweC+Z0A3rA80Cius1rIzDCZvSk3BiZ9pC2/42+Xzzbid38ZVr0N4T1ybr
HDCvmgkx8y6Yh6GMyF7KT5vHsQDjetKQBQZR+b2UtLyhNm91nzKuTutKlmSwEmhp
U/ApkJxV9dcI+XVcIhJgtEnRT4P6tA/Wb26s+bGM+fZCkTQ7c2XASH6bGt/jflIu
0+zNYN+H0BX/XZSROSSJchRY7bqVQSMB8Y9kmTpxshP1KY+DrbmRPREq1rfHuc4k
8GP7CfZuXY11ih5xDTaMPpBTUn6N52DZWjh04SLBr5zOISQ5rmL8cZqo//YDErgh
C1ZlMS0MyflFznWpeeBoaBX4s2DkyoD4hSaIAt/DXGw6ZSWIHfzzZHUQnPnbFtIJ
yPjaLidkkue4BEsyDo0//+ngI8ugn3ioZymFlP3SsfTwnmTECDuaioKV8pp1kiow
JpKzGsWYob157m2wpvxdd/H8Sy4W0Po/lha2LZmLlZ1BIcWY8kNk0gGbWJHLekej
IZgWZZmP7jcBhzW0eFJCJ5dtohIPN3+oSKgejx3Qt9zzwB8xJqGiPrgkzK4Us2bc
fqZ8DUoFFEuN5kdhT4r+fUBzow8pnz4hCSVWm3/2vOpCXHc7cn1bGUiDVVxEMJ4p
N7nC/J1MKaabTthbIHPp7SGDlrYF0fIq1+WxjhHwaR8vB0ErGOhw2lAxaPkcM7NR
Fnn431I/ofrd8f3oK+bFRCbG60t9XkG6A5cCXnGa6CkXf6feAuYbFdhNgo0/hsWx
aZexP0bXUcSVK0NcnIgrs/HuBZOILi/H9ubgOWTWcJG9peHZ5YTaAaRXOXljj9Kb
Bo41WUn8PxVJI2RgoV13Ko9aDmKc4kdTs9j5nbiUCNxfc1jNZ15xqO9fzkYx4M9C
XZQT/U5ieyU7nfWtfMBkc6O14coYB7zWDpQSXoKHDwn7ouZKnT0aGKaNNEKhtnpa
UBZKJ+2jL+kTI6WYiCeyECUggO3zMZIqRo7f2mW7i7vTV/cnUMXm9M8N3auI/SFF
UPIsdiO7IxRf6dyV8Mci6d0se7q93c4qAJGd4QbJXjANre5T0u2irMQEYL9abis+
iql+bxB+OB3fwhkw11deqTix8JviAXuLhJu5ndnJ+8fU8mj7Yf/1T8DamoKaiwgi
0Oa6fOwqnZ1snl9NfQJhRa30SA229HuJOjKqJ8qTzwmERn9V6BIY9NfZd/1quMDg
4sB2AwbRQdNyqhPZj98vukuIoOpbSCbbLy8868sel+vVJtYAD5POvFg7w+QRgfWH
znuWQx9UmWQfc6c09mbja2iQc3fX1sgFhEtKwdhAnyV1+HJufHyDtoPOsHkcRCZi
vIcxV0iHaRdOyVmm4ZEhZi9B2vVIClDoXpASGYFW5lUK5UW9wccG+bDcHa1h0m2Z
1KMO9gj+jLffxioOtjWauJPjSk1spUwdF9bNk2dnj4mUyFOGGMHtUSG+cNPxd+93
Uaf+pFcy9xB7BDIboihhi7deumrxVMTrxcb+xjMIFi51NpoNaDg5VzkC/b/sGLNh
M3IXhdl76ZRxzCRTcn0iwIym9GedZGJ0BD54fIVK+9XHGyJ9l8907I6/nUxtQ2MW
v2GnlDtp/QIo+rAZNF/TEjl/6aPJi9q3Gh5jBL12Ya204EaeOhFNWzerOaeZO/O7
H6Qmhi2diGKKOLzdQW0pl3pcX3ujG86xx2u4uvUOTqNXuFpd1AcmAsiBBq7WB5vK
9JtZ/kilRfEGZ4ct4b2y6+bXDoxr6j62T4UCu7/yyjdzi4qM8oKk3CXTcYHYw1xN
B3Ux2YPny2hhHE06Rv0DobmLGWGEeD0knHzCgRV4Z7WeDPJb9s79EjCTI/dy+fWn
kAu9/ffvKcepzjehV3Y6R3oWzJiLDFbYVGE0RPeCFLnYaB04aQnPYfkv76DsQC/b
RmqsORMoFrl3ejIM54ejzsemWKncXZlo0MxbBIKyhnbjR+RuniAcEFqk5xCLumc3
EjImSM+gNWS2GmaKvJZgK6dax+5f0rjW+LqtrJzkp46mqh8ZvBjpg/DQhXja55S+
d/laZIphqW+dSg/QK9Q3gIZkVB2N5oavw1vXyXGqkWwkmhznCPaPUM+wa4h2CvhQ
cNI2GAuzPIDGKhzhPD1nflL6Raa+0Y86EdQ40A5HZ9AEDprDM9l+13PJVqdt+EbU
Jxkc7qQabChDz7HVuS7ziHH01+ZfruQPVyOZlWr+wZJc7yyHrAb2C7q6eVQK2R9M
JoiKVdh3E6PBkxdLudrpdCtnrbjcdTI7WJN0HiruHu56LeI/cPC6oBbrZvVVADSc
42AxpsZC1mRR8zVplHAuqei82XQKsBQIbDj7YUwB7+A78TQuokoAGFCuzikLlWdh
fXnip/UFg0aQb3+6UjNL86AKw9mA7QZCRTQFsuYBsqp6xKcRbd8Kq0EXvVLWPChe
8yE/b/cPrhsyllPoz8XlZTaIW2380AF25BB0Ahu8emSTrteDG/vp+4NjC5SFt/4a
MGW6cfMnuO4kIUSH6QTgonE6SkxH4BjQsxLUYtevYGpLE+shGQscoq5CBq0w7rHd
I5+L9YPusEQJHGyfWOPER99Ksi2LArbJT8LAevwey3dnzvnsAkbhy+ioih2gClvx
cPZDjZtImQDQ9xaNAxYSYoQOp44epKfuDbgI03iHy2C8b4qB5L+9hQb0HBknShZt
qAVthxLL2X9kyu3/kyHxzcPgvTM8jg7Szal8NCFvmwghcVZecOw9aIfhI3OM+qG9
GKMnyevtSq260W7+jbClTbdsmyCFI/NVaVMnqMZKkpFwZoU73kbMvwCnSrLRxO+T
9Sur3Rp5n/IJ22eXfP28QG3Sq+zirFf59RB+Oxtpl+X7rUhZTKWoPNhAZWsaGLNb
OfDpl23TJXDYZ0Jfrcs/rVdvnQ6UZe67tRlDCzY0HOTxMVUhPE8Hd2JLAqrhyYC7
0+9/IjnPWPH/ST0B9MY7AbvNPJIhaXh80LyIobPUm2RTtlQ47Ew0IxPOqTnF8ZCT
+2+JfOaxOUo2U+OrbLNFIeqjG6NkeMDilmDF3s7ZvuDg1rnRuUTBoV0ddWABb/3Z
Y+c9YNJyqanNNAroZgAvxfXoqAhA5W7hkutgGo6WgmMEmOyLROPmOiaWxBrGoh5e
F/Cchgr1ummcioFGIY7OS1p7WvWV7E+9ft2v73wXpybi31XLsXnyz4hvUSRuUEpu
uy0NXCidKWe4jKADZfVSgOGLupwthXIMf9ldpf2wXujYyTufacwxMoMNGiRXNkG7
3u/3DynpqFPM6w4NdmWwgTPX3IBFlj7ngvdF/8oRVpn3mA+4btKZ+9/P7GNu+8oS
ox7Tlyu4LDICDzkntmMbwQjlAOg1/Nsz4AewotKmePPUYQKhsRXdMgeW8NYWFt+f
i4udOwVTj5OWrOxlTtIyP3V2HwO+gjvYvdjBow0gw+qiXLRB7EJEeofY6ep91zpk
3gUkbOEaNaYnXq0Up9tzFMlJp9VD37S/g0SzRqACs9s9uUq6EJ0PVIn1jIHfWpHG
htkJSe6jdVkHio55yqu45oEw3O/u7eyYYHzmw+NISYQeh9jRCDXNqS0AfTeYXrdm
19cfrFQTrEAcA0yn5Y6pdhKbPLoY9xfEeJcG4arNfYjh8WAvImFcmvz8H67lk5VF
NDJr9zJuHAC0iVMrh/WistZAhQiyy4jSgLpiJQzf46bqvmdjMt/9dI71o+oyi1Gv
5XVKyvaHimBbnz/kWdF/2LRXTvVafZ9F0vrA/t8fAV71BFMxZ1iWFwbzYmCS9H9z
iSK/Z5A3bc1SzZZo7UEE6vFA0SL77rC6ObebtZbUESRoNsWOO05u4IGldyLhpXdD
M34obPd2zYelBEp8AoZVWJm7V7h6zQE+Ndn8G7ulwJ+mJFfnm/M4UeLghRdlw5/r
AxBEFG0Qy8DSQpSJQ4nQyOd5qrk8LvZdvjULlhFMg/kJ1qXUtDrFsei1bSoLw92w
b8KGRrZcJf4BFdl0vvrscJitPmbXL7idDjIoEhKx7fRYGLr0wVTPA7f/PQtbJCF5
uxD053tZsfziyYpFtz6QMyvB4wX7MlkKootZPRDa72BRcnvb6pecGBsTMEP+zy+o
CE8vDa4xQYHp1zU6Adz1ZoFIT5C0qXUB4AKvdTRBc81Yy64x6NO441vewP3u0G/B
ajY7MnLfmqO0dhOON6VATxSgeiqQq1BiV+ai9/5wXxkQu6Xd8aTLRQmQo60agGe3
4SMjs0YoCWv+Ji4NsPoxsTz31WWVa71YqsYoZLAU1ysuzPOzm+vTyq9u0VCgiUCj
ihZY9TuF1JFqWLQBAFCGoMcglfCQIQk/nkIBCBaP4WbKRnLMeQb9x9qJDYbDT8QR
AJW8Pz3NNElfIQGW7pIMIySQ2vrYGt1pQmD+21fF9uNWS7H7400vdl7HVCjwxu5i
eUJjd+pmudAEr83gcU3ntpUh6EJJdbQ0MGPqBtUramEMGhWmX3Mxub9TP0gRmnbC
VJKBZu2IYGyAohdWi/+MqL7E2PZF93BmvopK9+ZHKFfNWjroz5qDkobDW/ry9I3E
Ab8wCq40h0AeGVj9tb7r6+qMe3UWt6xpxBrP3VX1alwP3F7Bvxz1iVkb0eAMXueG
ewnTWNXB00DmVgUu4Ockh+4fHIgTuIUF/aJ/ErcQ5iTB1oyVOP9r+iXalLhUhd/6
ufBru6fgNR30l0mNPN3K3EMpwQnIf8iNatsR0tIe/n4e6j5RdrhgnlFg1RLxTz5V
SGEk8C37BJqUfhb+M4HVG9PEsvp0+YH7KMEJMRkKkXPFfj9TH717x6oUh4zK3zZC
uhqEZ+OWKVqDzCnrjH00K89+HDQzyzGmUs14XKCIUqTpxCWhZuxQDThMcsdJKu7c
p533UMSBgHKNoNV95hBpAEWjlqhxhKOntKGcrCIUx1mIoPf2JmA58fT4oYHC1Tb8
N7WoAEXU+LofgRbVWgUxuc5V+d1EDu3prwOX3WQSaMd4rEJWgdHCAupfAHtAI6Xl
llBNM5BzoKeiafOzV69qJOq2eNKQLl/2gZwtceeLSiY+G9Tbq7HyXlnC8WYy+YVL
kXMGaUnsyTZ1ylTEsougwnEfTmxF+h2jBj2VoPhFg/Xp40cicD9Ihs0X259zW5/b
gUlPxtB6E8mgmRseCiGDLzAg60nmKL85y7Ql0MQckHVfdUrEJmgjfAUY0nIlzAfi
xrYJhs9o5o3vP14T/orFbqbHRAqmDZssaX4bDY16rhhPtUfM03D8qtIrn2t0aPad
ThcetT0RuEJrBgxSZhWpgsRob8/tw1p8HtPXhgq9DzIFXPPHU6St6SYC76AMfZFJ
AKKzxTrfT7yQQRYoo9CBngvMIAeRsZVLWLvuONH16eemEPxzcHnJgP+CVfow02/4
dPty9upPlRuF55VIdVbX9A4pk7ZwzoXzmCqp8nRCWxyQtch2n6JTFO7klBQ4fFnD
JWsDgTFOUVOZy01iHD4QwOY1EXylC/3VIR1M7knijXKgKanOkOTOF/NbMSBMaKvQ
JFGlkl885zjpaF6U3b9AdZ0bcrrjmXH0jaORgjBwVteR8NmlnRlVNvAp8+Pf2sZa
F8zi00CHjB7tDeNNY4y/xMJ565ODETizlV9PTIZ2IL+Yko9jNLIfxy8rouILtFRZ
idPWT8s3PbmTc8RLlxbkub4P1KUh2+8YOxJPCO4sRy59EhVbWhODQ6JRZcaQMRi9
2MOhrboBbzGep7kdwaZphGyxKxcU0Cqz+a1dKAxTfx37BvgITfp7M/wzJbDTmxfx
LOp6WQPXEJQGqv02ASWl67n0jn4Xy3U6SmELZ49TkNlpDWxbdOOW6a1rN2xxZ3vu
mXv014dL4CIvOx8KgaMeADQUIegPH578bCDxvfQq5mEY/aInuNnYpI0HZODigf7T
z9GltHJrsHYMUacJ+EnI7HxuYwtBppQsdvK9MP9Dj7i1OV6zhpy+ea6qh5ip8Uny
LQsscSaJs32+9V8e2sqDfS6wnKe/7+Yp5cV7yECZIwqgS/cO6RL2MjWnvECPcupp
XO6S5O9ivW3Dy9bbyVGPws5DWZ0dQ8Xztkr9GIV9RY/jxhsOWNVUCE+YZxbEVrAO
2Wai7ujhUwdnHUURajwZwrOSYKt0vjkAn56faXYeF4YzYE06/CnJiJYZeVNiZUn2
NS5bqVo6rYygGy7U0Nv7Q01F97gAl9LvzUfAqFWwdetpEAZmuR/RchdkG1ULmJf+
us9fzaFXxDoOd0XtBAy9oevakeI5+GYLjvgZet6Mvpj0z/kTGrz8MGG6RKmSnTFg
RmZh/TlN7Zp2eONibLZ2LwxztLmAH64rv4v8daZ33ddQ7RBOmHIlVMeiiznJGbxM
b3NGwRlZvLJM8jRfMfet8sojQdiBUfnXHYBM1+sCPzGUsWSahKJ0DJ9ah5jp+1FO
Vd3TLWzXDquC/Otv4svKTGT3LbNiQu44g0xFxVFf6hAgTDtCcCkzF4OBzVcbztUk
EVTO45taVvPgd939twDjlRed8M+MJzjGeVuuOmzq5G0nSpBp5rpfF/Z83qZ1bbpf
4vRN6LNo8eZ+naUSgST9ujLymNApH4n/HvOe6WvxT4ZibqIsWvgh9fF0WuAGF0Fj
Y10orEhRzBFupUuyS675ygkyI0rqWHQzfydmTxmA3Y65UEFCYwlZ1BrgUJlVv5gp
6rdfyJm8obY1O524RwV6QavCqWkTV2lneKj3WKfVtFix4QRGmG/rI0NCdksm6+Da
YW0CBo3e7fTgltKQOUeDsQGwQDoU+dchJMln2uVJBNxer1HHPj+Be+1yfBMj/Juv
+HlyFo/NPxoucAYEpTFr+42sHpm2njkANg3qkNZpsvAzR87Xp8+7309FQXU6kNx+
rpfJqe9y+oimboGlu8Z7O0g3HMB3DOF9e+W9GhFM9AKKl1F+jBqOv89DJkfBxIUq
u8iZ4mE2dp4gLRbvwPWFlhLhBdkwwGTHywsolK0pGf1hxx5E30baVsgn9vA1sTgz
BbHye31+IRAfVAT01eMzauWjwKWxvv2xgFBsQN1H85+a6/JEIkzS6m6ebn5hjrbA
e2CrSx8rcmrSzqE5QUP2VRKdFnKhksIGjIk8BbxpP21hiASk4GgiemANQosmX+7S
aJz73ajkWSzb4RAfD10DUS0m+i4GjXAFcZsMbC1HtAqqlRp6HmW1e1wiKl5TeYLe
B+s5RD8TBtQt2Si3+fqRlktmsVAQxa1O1XpjQukoaMjcDH9y3mjYRJ5d4R9C1iGp
/SY4ogj3L6wL8wBph5h2zrKAymYeVTD5cOTGs+2UlVWdqQMH2bvHaJwfX9Hq3G/N
glKyh40Rjm1j+sYUX7BgtnwVvraw/zVe5zIQMIEdBODXdlFxL2EINwl8AcBV1P0T
PxmzEF7vJUVG29q7b0N2FtJpQ8gj48PlLsxEwHUtQ6OLgVUaWDfz2qqMfrqXVwiP
+6SoSJLaoiLf3ewUFRt51W9FnbbmAi4qNkZBLhs7urv30YbPwrJCQsPRM60ktcRM
FbPu647lV/wA05pp9EClgL0aa5utOvcMbOBPUHp7WzJE4SxdhJdWwqfvCdpVdr1o
JuR8wGAOQ8wcDfFvtl/fuoJ9eJ6c52S0KKlY17t++MkUilf0mcJa5hwIpFz0Ppx2
eZWQyzIGAkvbXfoyNKoVX0PRmzztg1b7160UNYTQKhVFX84F92bxKJakthI1Ayc1
iePQ6Kcc6g3HggCPz3w1MzH0E/suhgC28+nThqyLxF08tRMEUij4VIOOHuHCDIek
/Ax0o0abtkattKm6uu2MPYSJsm+FF1OSQIxSqxKf3UXY9KTTrpyulLUyUEtEkPKs
Y/sfrVtqP2uhkEDzSbrNF71+Cq8AvSf/9XdBQumofpHHVN8f5yzlo4GjeqcXQhtD
7O3jxClOJuyDNC5gI7CWDWv2w+MFjVf9x7hCcjMfbmA=
`pragma protect end_protected
