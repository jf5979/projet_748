// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:04:25 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U1ihJVz3jJs6LtDJuk3/O8GjLOu0o6gMyfl3xv6CmmOZQiCJwXGVM8D0jD8bJNrd
JIXxEubvEZ88QhA8DC6GXbtKENzR7LzzQn/En0QZLBI8wZnpCDWDQQFx1l5CEAgN
BYBrxOqx8tY01KN82yzzz1JPZowaTnF/PxZGFBSJW3E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13840)
OsfE49tBd/Yr2L5uusKw8dsssg7LpffrbqQ0Fo9bRozGSlSYt7PNMsEOWx+EHLwC
HkzRiG4dVi2jCZlB+mJYM0A8B5YBkBhKSkFnvTMrMvfscajUmLxPv51bCs48a6CY
PtJuJV/P3OAC2TN5xPqGBhTLcpvTa/hg6QVVqTbwNibsqMxZLkDyr9XnLRZbHCbH
UnU8SRQ6d0k3/GGhBzuf6S3PPmEDGyE3DXNj+Gxrvva1Hultb6e3QKDK21CAHU9d
AQUO+H0KHnu2ochxVJEhur4xqZ7LNiKbbWu05ViBTH4S8Lj6wskimRjR8WZrBkGP
Lbhl5rg2YdVVg4SqFFavAgRIX5mTUo7wNvi+GfhU8+InQ91x3YRVZqwlHLDOllmV
fAJiDSNN3nOs+QFu74o7s8tkIYI0Epyq7Mh2pqPr2WSdaS+VXRI7v6GwFLMGQdY6
tZ5OIkb+Iw4ZhfVsVP7WD3SPqvOPtlnQJkwFpC4qBc8LhXFCRAxwQmXvjDtSnZtc
hpw6axK0rSIK1eEquCz+8hN1+oPU+sNHa4u6Mjz+6gczLB3P7ZywjLnzEPdXYPPm
jk/ojgIsxHG/hzvulyra5mBKJJKoYyKCJeO+ZelrTVUqe3TT1i32m0ISPS5RqcLd
3g/M/jYQLaMftEcpn7Fu44uYntChYhye4T1wtf2fmzyE8WaEr56uXPnM7Zx403+W
TzE1SQ0kMyNaybi66nRGB/IvmXEjbkvg3j2icc+fW0yqrKaeD3LQ5ztSZA5CdRFU
MplcbDpcnl2mD8uTHpK9KjHXgNcDTHRlNcTP7i28FMxjMerWwCCvbXs3edPB3njP
vzg+tKyDVyZXFqO0+iPVaddlCXkQxfLWUUccAHGIIGJXgS6l6vjsMw6Jb+ofo4Ss
m+I5uxWUdmMuzBHBFXWzowq4HL142nL800qDvsAKu7oQRyfJPLb8ZUZh8bOna4zN
I0uPW4B3yWB5/6BRSBwbsluAkB9ZpwXBs02YYV5jV9TNHBqIvWVkFvjuOQ56WjL+
L3lyH4Xa/JoFq2whUm45ZJcW2hdyda2zL+fcW7+aPrys9bI0TwwvBAsckXy62ILt
nlfpJHx2JqnHZB/IOREM5229lAlXwSZXmxfOZri98/EpU9AKUXhVy8VxRJm75gtn
JxS6WXUvlnz2Cv3tBRcESuCijDa3OqZ/qmuxDdev6jWWvb5DR6o4Ei8i1oBmR4bj
IVgiAUXRvq/pDy8FnJTw3X6nkSFLP/WbYl0XUbiGJ7NIkd9RH/mrsXT5kWg16UWd
vVudo42DVYvIdsoGVLdK2cCTUUCH3qVznxGYdK53W9k8FKVJ+3jX/Fw+lE+n5CcH
0Sbwmy6v7MagXTEZUlCvGGROsBePSpOx3oYcEgVUq2wH0El3P9dmhzzFWmjFSSji
zztxUfSUBCAMH1hKK1mVWZlWO5wyHjGbZyE6AwKC6CQJeygt1L0gAvaHhWfNLWKw
L+GXc4oMgxH3S+2RkrLP5rMoijXpyp5kozrkqBeE6wgLr7Y5CDSgfiaL9eiktpCN
M1x84E4U25COMmwPjRjSNw2oa1Hh2ivwqfmWNU8LGHHaZ4l1/aERWmVTA7PHbBBZ
ivl0j1wQ+pIBKladew2ipRXAzGMTfb9yKv8nSZ01wA9QUZcU5kMPn/SxbmSgEA6Q
4BSlhmIY8IT5s09w3m1/lxyxs+CxmvZbsGtTj4ohNCwj1d06PMTIqG1PjD7OwU4m
6iqvH6XY8ZCTCIVJ3Ld/AY7G/ohkarV8Z5kbEDe6Hvsdkg+mIU6whuwlJJd8dPDy
r/qzbeZlJYnB4g6PE07KlzyneQWk1z4oyfF6y5aEEEV/ac+PYV01r7AqlMQ3AUMH
SsmY+0bedgOjxFTGH9wE1BqU2A0vYR/Q6eUXdF/qusmiH+WVAyF6HKrwt2MW6qZ9
y1i0Q2QRC2IRuVgxl7RzS7t9Om1+/WPan1qCzf6pSnKBSawcTeDMKbor2DtZsDYl
K9/9w5KLJ3Uq7lw5+PPWQh8LssakIoCv/G85qhvt8O9E2hmHePPef56WLLtkpKEM
rXFRr8kPs+uJ24FNdD0o/6oy7lJEND9OI1HV0keDPzUkLt/qZpmzEzaogFJHZils
wHJBsZVFiuwtJqC1HB2GO2OcXKyqf8wuPW7EPm4V9avCaQlfr/Pr40fJ6bRT3m1b
iV4FglRTeJhMqGHkFv3INpWzU/wur48/+nS6Jk6jS5sObrUkY3ejF5n59P1hK0CG
HCeVsR7XnRqF4czZDVtY5axv9ANV5Gy+W+TEGr4OWQsRLD+vPuUs4zJKXUkvDMTn
v4e/M2HoY/6SG67ZJ71oTX1HAqt3FniaYehVVBwVCteZ/adetkV5qUW+N0f+yawE
tW4zkoniprOIqK7vK2Gysi9Hzu5ewpMhOddPKpAM2FtTaGAPKdpTxopy8r7DOOBy
lu+iVQniNRsZcM0DNNDtepvqBegpm3BBqDdYUbCetqxGxVLnr5hukzEgKeB1WloN
ypJL8MYK3ZyHm59y5XSD7fr+Qa17OOXWyXfXzwgOyqS6lOdHSG2Ydpz2rKhe4j11
YKvUedgnvPIyt9QBo+2NEeB89B4CYBUydBhpueRQHVVgtUeTANhES+QbyKYu2hW0
cYSB1GjFGyf3/MNdcbR4RVWcwEvOc4lkSdfF3u4ISc6ESL31DEK7gdlujtszV9/Q
pviucgKK0dGJVC/+mppmNWczXBFZ13H5mxEkXH1B0mQ0JhpPoVZBcjOyfC1PCRZy
BXIBoxFcHe4IQVJnBXvKDlc/kzeJRaz7Z0si7PsU56dISoNwK0ra+nmFVOLjjln0
F5TYfb82+PAy2qbDMpVd8P7Bn8KzhI3JzgrjAzjKCqOLtNXmEfdV5RC5w/QYMe1U
4dJlykhZSLkpci9W5rXTHtKUAVreND7B4Fi8MISBnpO2Bo8dhbY50/vs/5Gk/m4U
9pwwxSIMWiQ5zNsxccDG0GcwPhsr7E1Cx9EaGbBKtN6cLdHPcz5ilxZBno9oND9y
eSyoyc0SzRsJtFAIiIARG9drlOPSG/5VVt74AHt1Ff6BmCI1Osd8ojLEa398xBsm
dZzqvfQdgY8IWgjfe0uf58l7uFBsXcAyqY+7P8Vp1gIHftnJmkcat8b28t7kBTrL
jXI1rJWknNv8h/f3uWI9aHejXHJsAyoWIvBPVWoNFnYxUWVOMq8XlR6cPPeUD7hb
lkz2N8kpF0EMdgEBAcrA+ry45IKuRsxgNiqITqtsXCyrYFk9y4vifelJyqqo++WI
h+GKQJMczdXFFYPgGKXFtnDAn7YIWp3NsJ6s/ppbh9EYyFpjno3gie/w8sC0B9hK
TWZ6uW1AUsxE8rnjxpEtuwlEkXgJ0OWqLkF/Zo3L4/PdutUWZU6K6Dr2tYR3WCJy
LiDPe0jH4OpkWJ5AVILJJfi6CwVNzwlCHu5RgH20y5ADxg18VRgIT8I1B70Env1b
1DECPyvFEYZ4HyFqHWU4x8WKxtE6fcR+ae2gDcI/fFwgj7vbk4szD/6eh2Mq1Ix5
6yRTsrnAK0Qee00JmPd7jY5HhqtIz3xPWH4gFd8j6FwpJhQ4QOFq+ZiYJNf73Sxu
lIlgut1SfDy1L25VN2g0fdmSjUfQx0w5KltlXhg16IfdPPDNtA4ImyYqnDYhee40
P0t5i4H5jSZjL9wL45le2LoJ9b9F7el6OPirUtiO8AmBJ9J4HniFDXzPkrITxwVK
Wl/sz2HtaS/YYKKxQ6VPhZwUrgb1KtUQznREbCttqvQH9JKsijuU7UHQrlBlQTmb
K9PXrwgJD8iAkSbmIqy7rmJSsoPUoHKLe+ZAcOBctRGcmFvxC3uS3KP8NKnRKEad
sxzwuZb4w+x5ksAtATXCAnMYGioztTYLV/4MVlQqZFVpXUVFsgfrU1r4Q6Uei1bH
1SFpjWUPnoS3mTNAkn1eMsExRhP2byGfo1RK8H41ERGPl5fzhITC/WZfyHDBdyu/
iMwpvJI8Khrdqr3X4pnfoKfyxdfDO+6zSqt6+O/Zj1m+SWd3gRIsRDqrdCCWVl/c
BI35r+OEVhHU5ychoTxxG3AK5o1Qb4B0IfSalk1Pa4u2zf7xIl9bqy9epPPYBBx1
CbgMZGEBmHRfWI6jqxgYnoqT10S/xwrJL0KK7XNKheW7Wqkvz7orlleqzFVHjWvg
EaI+OmATcBSWFfHqqU6XH5KL+oTLjuLFGtN449L3K2zx2WPO6poeRCvt1VkZxdF8
/dvNOCpqQupaerzjIrQgA1GIOe/ERl+8rvhUtpKf0AKutDWqztsW12b2pb72FWnB
OuqyeaBmjcfy8WCeMiR0sfbElIxkea9HnYsqBhxUTmdxRtQOpmU7spKuH+4E7GZH
DWgv+NosMTK9T9KBmIPF9tJemDF0fb7GOCDefyGG0BJFlLZLIFCxpgxPXiw/jjvv
mVcCVRVj3a86tRhlIUXGqitLFmfrkXtNuNAq75c6SzktV4d3hr62Jf+YowDJC86+
uIE9R329MB1RLAFQDT1dbr0JGeNWOWgV4Pv42eKUDtZ4VeAQwVmiOr9c9fVcPnyM
eIiYXlV3ICkMPR1S7WELlAbaaV1WCT30n59aKJRSxxMS46rTPAhtgFLA0YaeHYaa
Y62AbAHbjrBXKVOPIC1umoxAJdx1JPAAjwH+pEP4MUBGWctHybW9MsqwbUnlpAen
Lhm9U4YvAEqX1iq+8AIqGB9pUtsRlEEv/OeLiJ5ej46DOzHUr3WAqmkYnO4UrpBy
gwkA27NXB6bhJpa7CgnhyssuuYRmuZD+utcdHCpczsvBUBUGkmI8VNgZ5xilWWH9
mbJQIcxlS1DyiA23/U+GClwizFMZSrVVhulccHAYCmv2xx1wPLKJyBgA0nzNVqu7
RU1PrvTxxZSjW5h2vuMhOrHNJSIUST+8D5/27ptOPq2D0bEAM3W6ch60uWohdQqm
t+C0taRIkvZAlEjK/A/E5f9Z0fIzl2k2icwJw60tvUFDbg1Ft1zmw2a9419YSN/T
DcbVdJBvyagioV/3WlxIENjH9aP+EoRymhN1rwl/rO1hR2VMrQfGY2lpIfYBMOFh
3IgCOX85wsDT4tBi0nP9sgvyEMp0uwt+Evxxp1oGdre73hRP7yxuUypvkdkDaoDR
sAnIKBUcTpBLJiEETXFVEyQuw7GxwN2ESbgK0N2V0ZaUhvFWZ20snIbooJFTz8o/
ro6L3EsCtuuIQftHV87QEnGoMBQyqSdq3v2EZNXTK0ysyD4r7jv6fNvwE/m3VGOG
zkGPm6nJkyraMoF1mQ6qx/WuPaDgh1ji6KNFjvb/YEk+8RwCwF1fj3wYt881FLTM
HntI73xO/BsmtLO9bWw9Q0bhIJG18VwQwaPKbiPRK0K0x8ZdPzElVQV1uh9RucXM
tXmpCEEo3/kkyoHUaaIDcHRcwK9PnKc+rVVDV2H6mwrKWFq3w5yRsHd9Gc9o6QI6
S8wgqyy3Q4I8EMrEsuFNGTZgGr3S+cG4OzUczxenoBBLJ46te4hAVG3IQ8Mj4J8h
MI6ZYgNpW0qfo3uPhMzyErWYS+ZrCMCFiY5yfUKturaypjQe+kAiWw8UEGOwmCyF
OawXaTjVsBrJ5iAaLw5Th4I2Rrr5ssEf7CAFJyd7bYuBaoRhyr4IlAG+ohaAvnzm
NYUs6mlOrFhm4F7lhAD8fcW8VdNeyLX3rYSel+1E/h9HQgrlvVMvBYSQzGB535Tf
Tl3aZN/62hwSPyTcqXyo/loglYkESGlqYsqdMaTv9+FHLTBaEilwrYot9dfCQSsT
C/Vab7EgdyeFxOpFVKE0pNCX44h907TxIUYPhwq6rKlXFttHsKfY2K0019OWe4vG
ULjCR7doTl/axPCNIIGX3jSpvgDzsHlvQU5Uw1zvEAe+r96mspa3gDhvPRkslJSV
IqRxNCLSVA1VyNAd3SjTpZSZOzptGRgO/XHmt3QRuL/RWvDIuEaiX0Jnmo9iTlkT
DkqR3hCKCXmuvg220IA0czbrmew/duXpFeUhgK3XSITtvcUC/D6QXwT9A9fNLztb
3u7s7aDqctfyGrM95lmvnBVATjivHbod25nhCJlXeFmtPmHQDmmqWLBYWVN7ABV7
gmsSPN6y9Y6EOgG8U/XdgMeWPrQtyddIyGr+AqD4Yb3XH59Cbue4cUNbdpI+FZlj
TPibeHR+aFOqE72rYQhmCLBBMY0RGlHzRsLgRvWUuRcezmmVb7vpkRXaulGYjsgY
kEl3kkFPoi1gHy4Xl2fW1LYgk/tUFqVFoI7Ryf3weyYA4xzCCY0NF4pV/ivqAWB2
wdqPMM5KSFHiGlyQX8woTA28wWc1Mu3NzvPbtDLwXl/VnLy02EXU9C1SLLcyXp2C
wxTqP135n+BWa3H9QtbW3gPF+ILxPeeZzbc0l6Ls4DMjqApJTkvrds+33ZUPNcCM
oxHUVbCITDlrdMxktoohEQ9z5ugFLB49rPKMyH4NfJ5HAvPpnumStSRGfpFRHd7D
OvXpiJ994oI5FA25nA0ZviZCgx7YqH590vcZS+2LJNM5Zmjq6oF9yAcbp2id/SDx
pP8d8eEIv+YxkHr7hCyWt26fVG6QagHAy2+XF7UyJzdZ+Udl3XYKbTM6iJQNGBVi
ZE+WyENYsb0hPiaMwtCjoLnYYr+u572Szyb7WtuQwDRft4O2YiF2JswWrWQgYNvD
FBf2Ru6FZalPivlzvR0MxiY76JH0AfodPH6fGsM1/9k9pL6TWQ0Lpr17KkzYM/0e
CfD1yYCUZN1a5Zj8JFBW14qBYN3RupfRisvkGhrKbiekIHT4LbxOwWuoUWrCJheQ
cdDMzxmmMkaOMp2ezq4vPrdndy8opYR6QDQdXuLOp3L5+EyJO/ffCAYGJG07ZPdh
XQrbimUr0cq5SV0wGX99Xds+uuOXvORm117yweshrCOhAs+opYQCopQJU7+Nxgeo
H1RhFZCXr40TbMQpzHHQOs+9zu/6BsaWji9wpdgwrYLWQYjagI92EZHrCrZt8gpI
r1rpQzJFZufGTyxjpy01d4sdTSulqowV6VGNUWlfJy44JqofxFYnXZOxEE+s2OXP
8+5Egsl+FEapT9vApXMZkP/eXViBeVrhLhi870bKcpYTFFvqLWcbLXbNKi40hXFh
IuHMw/qzEQ8Zv4w5aMcsRpBKDgvGhr11JIjUKU+lBOK8j794Xpd83+5j3Td31mmH
POYe4djCHf4pawZvBf98hY27GzwnQcR4QAfDEOfG6QRS3L0aqloMhVTWU/aFeKFN
0plaNJesN4sYgl2hzHU2AcvRlYrSGGoMOZMQSxG59QrZ/dAsnHx+EqLrHSutp2/i
fsmXl4rx7S9a/yrn5ywOXiZGEaUz6xHtX+hUx1vVNdVawu6pGohTeyK32UbhskSu
6RVYvvfg3bdRK1PrFpg1EufystMi665M0Htafr48vVZVl6L3a6a4hhzNlr/OMDUg
PhKzu0nZT65ZxVzYGlpa0WeLau32uM0OptfaVRy5upsDBSui9aniH6xUgY4UCOE+
6B7Hy1MtwhJxleYXZv79koFzz674K3sJSHo8wgE/RLz4AspjrWlFle/yvLR+gsb2
KAisbUv6vdSPnQPJP0sqSD3I+M3AdzdjzXXkB9dPJcVk+ZhHKj6vB53f3JUzjtYR
6uGDanQFjrMR1Lxm9utMZRGI2MwjTZMbJe/KE9h4YGHYIyZ4GJKFwhCpgCy4YsvZ
/0EWLghZLAjuKHHGqvCVqCSc+ehqqMJ/vGq4G4EI8SZFfwHb4lJ2Zupd8DLAr2gV
OSd+KGcnXSWY6AiXFtuRVt77pduBYgT7v37QbXFzS76HKgURpXCBO7hgt+kcYk7u
DVLZ/MR8VWzSoTRYg2WdtD+JuqJkk3Wy8fMYa+5KLDmqiH3FMWGleblOmxG00DC7
ZXcQ7mwi5o4ZTqz18YwRYkdina4wvnW7hT0nMdhJDJb0YymseYyzRXImUbNb4lEZ
cVO7Y7v5D3Spje9YfgZrQSK01wyerToCKt+JnnPlVUOF7QlsabXbvZRYreWbmWnv
2caILbee625TuqDgYGQBhPiSrIJHPEaC5wxvZRQNfWKyD3+pa1TZ0+ds/dBMW42k
jKPTI2rAswrn1Mf/ksHeTdQ5iAoh8sO8zZYn33QhhmCk77eSIZRKqM18WAK9VqdR
IOeyqikmCbgcyAgIVDMMEtH/deifTeihV2BojQom3GvJP/HBe4lIGdD5La2xfS1J
C+psRsOR7NXssJRKdwCQudwu580e2mYlzpnZ8pCNFdUXIgioRTzdYUVU/242GSdl
DwNPt6YX1yaeddXNRLHTMNSQuM3z7qsfg/zOmsnILeG8iv1IIoadOoaaIZ89gr8d
fNnZde4IvZi+NFwuvFUOHkOaSiTPLiIcYfLMHAur+SsY0s3cMqo2aMMKEOC77vVC
AvM87nc9vGnL57GOK8zm3gsBa9IurC/F3uxYuWU/2N4nXTG8ICp5EwU2BLnlm1cI
GqeoIdyofm/pWBSzDO4/dRFkG3hZwSM4iyYD2RHD+dlVUfhjY3QE+K4/nHSyRGgi
cLvA+qkNC1EOK1nU57O4XXzs8oZEuH91ZzOjFGhhcMMV5kBrLMuudDDnLNR5mKI0
FPZYNYdPmhUgAUe3/xk3v+jTgxGd7+rUPV/v5ABmU4imI6wW6h8DIqoWqTc4HMdD
Ja2R7RBFvXNYLSjQ5r2xLgL2OAOata7AZiCY0vi+qpXd9scg1swFJoOmY9zqYF63
uYve5ltoHrk0VJ21ANaEYC72uVRaSBitK4avyD0LyjVJCGOse9yfHcfgwAzcWbjw
WEtNJKmPuQ3XV0uVGmiMrCPr31tiGhmnlSdUnQKEiiqL+3xQnMraCZ23puiSR2e6
f44H5QvSbOC43G6zOzecknm8Y8e5OPAxNvdUW9OkQU/kBcv+BTVe6gTsnUMfpLQ7
yz63ao3rhfUn0v+bcBzNcwTcrd31jSO1qgQo1C5P1Z9Qal+W+6qu4j7D8Wdrtsxq
mzhRl7QCB+rA23oQxstQ1bGVYy8wyv7B9pdmN6aYUWz33qzWyNoXyUh/WzE+TkPI
n3z0ERiHAR1jYU1Yj2INFIr3Am36gS9gtHZTWODOwZDjEmUWuKe608p7XETE2u+q
vsXZBgIlWX1ec2brEVBKtqeViG6jzOhuzkMZnds7IGhl+yW6jJmO5I963rsd1KYq
/yMkK+WrSE/keZKIPMumOXQtXi7cROTWdh0EIwLrd6e4+T92v3VtPUikx6g+H9fz
bmEP3icsqGaKE/VrqE47GDJv8DC/Z564ScuyenpuT6luJEo1TDCR39wVtPpDb+ac
i1uOtwl6Xt8UuK/uoFUKwWGZ+SToQjrhguQYVNtibHLgs2bbBJu2b6OqTxada0GV
XG2YP8KH4INPIIFCIUI+xA4vhFU3zB/fdhUHd45LTNaXKo2jRDfpSpEECmfRS016
Cfb6yF7zxdM5+nk8J0xrzEjhkQUllbrw8YK7bW6fMFWgnd6/p4WvnHhB+eY6rXYE
qbqMYTY6RfZCUDB+ERBudi7kg9ktOFmVhTVyfCRrT8thvvlIw4V6NscIY7wlB8+V
XJz4WFeKLd/hPSv06Zb4/p5dh8Xc3jbWEI9D2Hz+qBzUPowrVsETGsVn2BnQmSGd
23o8iz8AKlILfl0EmiCHXqrF2R3LMJJYZT9Ks6wNR7gFjmjj/UAZaZyP7D3s+ZRl
v1OCoR5MY2BgowXjsS2UME2roNIHQmnuvQ+SvDh+M5wxmZxYMiTgr5vnH/Krvvl5
g876gQm43nslqEOhfGa9CnxQDIFiqKaw5hO7nXQWgz6G3NoAsjAtPa4+tzBZ0x0w
qmqNarx/qy85+MEPLhQ7D+X5zOvtP9LSdj/54giyXmbAQ4KNOXtE8oZfdO0tcXZV
dLF0/BxtLKpyRXU4yUSLUCys8KAF25/mEJwQnto/9dgD9k5/3VWWy7rBCLYWJtTK
ngPLqRJpL4bAbbohYgWoUFjNujS+kR8lI3srjUEWz6nd3bu6sPwpjDnzNPm8Ehga
ia27lxx5qCg6RSCR8edD/dwyI8+CTCurKnZ/zP1vP862UBjfQGESWxT5zT4N2uOP
UBsAWheK7jyOtqUIGxz2V9u2vnh+T4BRwsFsgiMJzUpMOsZPC+eNyBNY0zlgQhp/
CI9dD/3kEYFEOWIUei3NfF7P8lZ+aQPS1v5hI00nBMZKC6+4C+NnPfPvAJbw6/M0
myduns8yUCfdckX69WL8Z58NbWbJEPIkc+x9S9vD/1AuypQcRckcy/C1CJ2nMUGP
gfnuMqpuWCnd3dtUvO8U+NVUlqwlclrCJ13NdPF7yNp95FQIsNV+dTWC393JgUyz
r1qlYU4Ej+I3HG0d+upQObfQB9fhsP0kx4Shm4G3c6A9FkmFq1lfrPel/9vLRRuN
LcnXOZ649MLwYTRlvhdu9QWIylH29Z4lIeFH5Q4+/WAhPiUrPK2Mji6cqDX3abr7
YjV7WH0ZKdsOWzKqVfodLpgpnWMD0bJsiTcICfbIPlJbLlk4J52YjPzwxcO1lcAL
jquQHu2eNENRvJSgZt1MGuh1s5Izry0mMd8YQbhr1NyvawdpkZkPktwr1qkVU7Nd
VMu8SzSBodjT3jBrgSbdMCX0nbG9U7POmb/SzEw9be+22vCXDt79AzhmMIKLLAA6
u8G+ihXHJ1imLlp+219em7GMPoRNjjFu0RSfqgZHP6mL5ba/HmMZdHhD7rna42K8
jCLKff9IRwFLzneVI87mvTCjjZfoo+/aoeX8B5887vRUH4qtr6QArOBj52E3wlfs
s61JanFDDDaJQiG3vi+tE+NCTKX/VdF00NeKEEaqNXSnl0iVkVI0gVnOMatZ3PzK
eAoyxQCpH1KfzhqlNnIsI0uTnPEkWKGydYvGBemRVFbiV2TYML7GZcsRayKWNh8T
gmlxl5Gf1DnNldTbEkK9CTSd2c6BEGyMqfTK0mDuOxGsklEri8wdUhJha8u55Am0
g+Q64O5DBv/uhcEvBfmGVkWsdGfvpPMpeZEPWhs56LkH30t3wphpTO1SNKHguno0
LkWBIaz5WQtMk/ysqT8JuPm0NtbOMn7xmIDGRNgcQHEZ5uCJ+6NmE19kGm6AOQBa
9fJ4S+1KRpbcLB4RTDB6hG+y/Aq9HwQsaXwnAjeMyOyjpUTS7vwlJl2EfpuD6jaQ
HKr84cOBF+Ayi9adypT7xxXqygr2LeMPoeCYXQmAPyeH+l+piMl3UdgrujlXHTMG
IM3pvu6kIoISUrjgpP6h3etMK3fFNISt+7ggRLyir74OqDODyIvZIw8zT56mFjvw
7aETGvIeP1XBTfEyitrQ2EHmffTdkD8CGfoMDYgIWrliVB6nKkExsCAS3WqTHMva
YGsFepvF4qNqkLXMViZRx3cXZGjYie5HgiRzEXzonw0fgW9vXolyBOhBeNkq1TVa
75akJNZfDz3i9Q11Pc3pO20QuezXoG6u62JtUEME4WZrI7JGqOtcYvQhO0lLV3JZ
mRCPxjUBsYY0miu0JCLbLb+0chY/k5S+vGtGrUkGF/luAu21Gtpmq5Sa/CydVzMO
Q/ImZio47kNiX2OYcvoThRj3o+omzqYgDkn3/lvjxHf7FMM4HVJYvkzANs1+2LLy
5a4lV6pT2FUBvB8yX4VtlC0tzf6ArA6uC6uhtErOWf5SngqA5Dj8CfnRvXSOaOg3
ao35Xjxqteen5UGqD9Pg4AzyLS29CWydaWDl1e/WvdBlBE8n3wyTBoI2on6V+1HJ
WmGLfpv/Z9heUE2HH1CTBWk5/RLRMoSZnMexAixhEYCqA4KOrHjCLnZOTjOGGAzy
MQalIIko8MHqj1ylGfNwtaUpZieMAANGHwiznpQ1Fy4DAJbBkenVqrO3IhtGoYKl
wlf1DQVx9BBSnK0Im/w5zDGefV+LFdh/8YCe7QSSTH6fEMOvzeRfrlNi7JJpTFWV
5syi1IjBfFX6DGrzraG1TV+7b6Mkln+feaSiHhqbxcNMMPxiF4MAwtU5VnsDvGbC
yi3pVNhg0e1BDZWpDhAeQlgocQpSTanF4LwHrV8eko/9a2JSOfidFYknlquXwQ0w
senpNDHSMx6AyoOA3indI7GTrxRmSzy94NUHtPLzK1lpuvqrb49sxG+TSfxgh2r4
untTLLJjawKwUtR31t/jcqFU2gIn3rKIXcE+mZDLQ91XBcdI8IOYRP/YBfYwGt3a
uMrCPWvoIS81X+SmXX2X2k+nNEfUrca5uDqbgWwS7St0d1h0UVa87F0SLQAPhsPi
T5fbhbwUJFlsZOXoOfuNIOG2BVngGFp0V2bblZlZyeH5iJUhCDI+DaIVma7TU1Iu
sUHeGxx6Ayz/QwJjVdWbHgMnVrFFP+I6o2d62noHZbAlLwKj6Ckn/YRtHzK9R4mC
EStJOxEx874uZfP4Tkq/htoduCrT6WFHGh2MrIF/78/+RPTTKwmlS+lG1aQptO9Z
savz1n5NhgXX0NEtJBx5qB9AThJ3eLPmPoPZcEJFMrgygY1cyo70f50xlR96/vM+
FuQSm173xiOtGyjqt/OMZALoi/sC3SjklFTrzx2McnsBDC+Fd/1kz6IFkAZukMQW
NZdzcIIpC9+YJYQ4fwENuJBqvzQ/bzX70vYfKcjbNn7QhueAw9XmJQH6Vl9FFr3U
a+GXH7OGSBAaBOePLRWyAvza6KZe/Jx+ruHMa+xfF0VsgOKa9dxFO3mY7R/Kvbl0
UBrERTvrs9GzTqE+lbvB0HjCienee+/8nVZID+WgrZbDJC0QPytOFGrAIlOa0i/c
NZYe39/DyR++W6oW3v22S3IeYY3Fl0nZj2Xr4SFzOQksdvmbnpTmwSHQAPXBIYpM
LGe2W8E9idc+rvUWpWlU9EUY/pLWIqt5KSCliroZcftaMgIV/8UH8fytrfmZPPbz
FxCWHePthMFN23XFJvqm23yVPn8ymqBeQ8KsLxhF09GV/UxpCfPxhVV//my/ds+b
XWQf1KQQDnF2L+DjAY5RMQlLzDYkdLrR2KJ/TrboUFMFrICY6g4p/a7O+9S1fX0q
OFk9lcg4dUJsPsmZE+gvI+JUirHVlEHYNmno96aLsz1yktx49mDNBpjAqzSxPg8Z
iG4sjaRM4j5Nm0Ex2sZQpIj9stUz50nCZtBtKydZwxd6R+UTj/bSImBeif9fmVUK
ydek346HxZngIDKl3BP9LZ0DH1xQAF8SQT+DWkBvdio3FvOmI9tWDZWp0LDfrgxb
BzrWsjAOXgOYEqnLR0Y7YEqMPAmNssujXIgtNrChuCnTyL5g224HCPqhr4lPX8l5
GaG0n33Nyhc1djYY/ki1NTmTf9Gyn8mnik9/i0XZm8m25LMDn5cb2z91A+uYNaIW
sdw8f1bYvF/4J2tptd7L+8v8JoMGGt44nl62WZeqPMszPgh57jVd22ARnfhMeuFJ
QvP/itY6EAwd20e8tePDxC3I3PgOJHN4yAV2d8xvQY+2d9Ii1GR6wVTk7cPnRpPn
wFbl6h3CgObAQdix36sBsQtRz/arUgWc38QzaSUJnJA3nUWHYMYJiqhWqoLWbb3R
TeF9s2DE3Z1KUPcMAu9an8Ua37UOM5One3tQcHE/8K/epEjzxcjSefGmoaOS0K+P
LVVlwDOsfodfRUdZfFRoMNih/4M23OrdSJFnln5Oc3PBCJx6m83qktj6lNErX+bv
mkTLfW+1tBQKRWxJxIwD6AOAcFyjKI7uDkr0w+d/nIWFVTHNU7DHiEM2MdFDI/1d
YewMcWGMEdgxnlLtr57S9zg9QX8dWNVoRFGgB/mtC6rctvDYQED1FKSwrXTEAEM/
Zrb/EDAbG2rNXbXVAGVs9If3cYyInQhlf4Nl3JYbRlwRkeqxmUh68n5LDavTApdQ
vp7Yaon5043mlo1PEL2GutmYyWf7lI77dUiBji5Xmh4t4S/OssJVv6wfF8QF0MG8
rTrO4FdAX2Q/wqJ/RUiLdrghIoHuy+GmBbA1X5DMnB0K2w1xH/fAAsz2lEx4AfQp
Ej7JJm0BXd0gfQTyl4zc8aHoHDKn9qh4Vz8gboTI0/vG/s6gAM+/ga2ADN8nYlw8
mryBAENR1ar00MRXmNiloghjhJm4y7ShU2tQ89CgzbYFYy5oCxr4BqDfdrTjj9tm
Rl5/SzmDYodzbbo+1YAjWXTdJMAceZRc/Xlcu7XV+hbzqnM4v7ea4ditbq3jszzy
I0x9xFBZI0gKOGXGeycj4r4DZuN+JbmP/w5CP2BtV2HrHT+4BhsORA6xAmUZbm/5
5kj+iVBF9fYe7QjV5jlfPrr8BcEDkv4eRy3+VjaUFb3MqsmO4Ev7Mikfw/bb/JbT
3U3KJ4dF76M8gj8rVOkwBb0YbicGQ4zdiqVpPD90zYAdiTYX1g9ehxydpyDPT0I9
pGBFaBGmYagoV5aIR72uy5E3jqepjxm/54muuhBH6U/1q7R6zjLjNSZtyvC5NKTa
NmyAP/G8FdN666S1MSEwpF3W1IWLxN/TnBNSMHc0dMEIZD4Vz8eGCbCRXHA/g9hy
1wgiE+A47cnh7fa//xDa+2KXCkEsvJBXDnD9MTTy9PouoOCu2Y55TZ/NiHemLhNZ
SGskw3utWD6teVdHIdNGCQWcBv0knlaQ1S2QSZe2Dlv8ykzOoWLdR7F+Lu2WUWH6
e/xkLJKnORw+GVqAdUeo+fimgLAMYAktsH++7zSk5/lPVhryJkOaOw07EfOGD9bD
5l6Ahik3V8c9LgbThNgtQHqD87RZ/A2nvIiAfG+Xc4fkisRHKG2fKlNqM9d3XUhx
khJszzGL/HXGqIafLj/+htRQ9IOp4I4dIEWS7161JCo4V8bVW+GFHQ52UnYFZFAN
r3KYaCWUkxMym2b0bGuNlbCeTTztqbYyJEMEk3h+m27+Nl7M05wsQ02NseCIh8qU
2cCEPhl347aPZYsldLoVu0/7AFPgGE6Fa++1KqeDcKPbG35yRlL5KUuASFbYQLJA
5OpvW8ptqgdMXjN0n0zzWWG0Z54BfMyscHsiMK13uMo79bFwTEq2e0ZCgdwRnUJD
PuN8ybTmBTM7T/iPfBDxjtQz7dYcMwTybuOb0OuWy1tKhoGXKaJM3CBxN0cd8cry
TOc+YLJ2tJPkPMA+BtL2faIALlGW2s5hw0jSst4VoMDU44IO5yWbQLQlHznzpdxB
htHsT8iFhat6LwzL1563QtKII97R1yozndK4KizR7NZEg7iBdHA6qIa7KpsfSohv
ejImBTUo10R5Mq2QQ0h3+sh02peTi+iLpErQLxCrsDUORpoecO4cJv8OTONKLwHf
KAhsz+HgFG6c0fp/RVPsbkaABYbGfw91Yvey/3Gco/e4ZR5FsHup08qrovQflwF4
uEytANuhwXgjU7C6zIn19W7x7n3euiqawu2c5Rha0EgIZhij7qSnp4+O92FYCXrw
zF/PrjTjFHLoFdsYzPfNRXm0dzcA4Iusez495wYG0kvVnfVejLaByneB/SHRV8ga
5GZ9clYrAR9MCi3+iD2nxovKmfp0DpmboHdgMRSSJ7jeN/9SsUEO/MmjfIVmUQ/3
of0c6rilC3P0oGFrpooX3IzHV1IeaVoFNPFONBLHGYRp0A73kRZtt9Lt6zykm4/h
q2kec1dOB9U4o9wXe5KSYfBOz11tgZzKhenlx+LlAcriUrKvHCMUR4fEXqRWjSFg
xU41cX3Epip2BAH1HSmOrcMeyR7bUKoNHfEK5BwYy3xleJ1ajFD3h7vi8y/9KtEg
6LkcBMebuH7ReiNkIP1/PjwHyXk7b9loXlACOmtirSaqSJ9i+cDQ7XX9Cm4T2fPT
o2dwQr6AJqlEjoil/STDJBY0HoQJFCNfR6HUGMp5giu0qC9u+5OfqoQSgsR0RY3y
FyXpHlR8vcbjkIzsDw2zIReW8S8Zk+6l3XY22duHaP0dj3bcKNMKi6YxDhc0qAfL
DAYSevsM2DVXhXQEY31ACmbZCaaOLhY9R9OccomwsgDN++MFjH26ezILZDOta+YZ
bK97Yrt61pydNJ9yFD0Fq6TqWFKjINuG22cqMKmyvs7T8BX3qO0GXtzE5EuLHyYp
LmkNOlI4EpoUMI8/lrkr6NIzQ0dG+dU31CPQJQiI4Q82KvdxdxUvsXamj14UHogB
SzbThCdZ8bIZnvH27djr75iU/P5/1zfeDi4aF8J18G8WvqqppF1vv3E+Rw36ppat
M4gd/6hC95cJIkWO/rtioWbOybOWsxyv59s4IyGqtGwW/6YrmFqdLNpAuJduFAxr
+1FHkEu4aghS0G0l18l1Yk4iwm1J/2WIWOv7YYN29uVeKAD5x56zobFqrS260dHm
IU4S1dp5EQKRw5LSxL5StfU2ASwsfkK9/673DM5CWGYXE9Gx9ELbSICZhJR+8eZK
w2MccphXryWn8C73nyjPLVObGXm3O0EQrv2ykuP4wD8U68BCozslgIpXqQmaWzzL
LyAhWYL3e8gXtay5VIt7gun5bsDYl3lO2/M0v0SMbyRpOYeRJju3Dxn732Xkivw/
Iyh0ekguG3VlDAtmY202OF3qIp0NCQ8eM1aG3HU9KewEJ3Vd1fRptGsZgKa8yh+u
jFVJ9BfLFF+qOjKoe/lEFEN0/hGqt92QMOKnq+qIYMkEhwWlz25p/FvHxopObRz/
YzXUMlmUxb5V0iRWjQlzaKf4KjkX++Yn5hPS2DfpIabTqMXD263dmJCLL9sRlKE8
2u1AYVLM9yHynZdm+8ByDXchDiMHE+U9chA6XsS1THDipPsSgfmVCuFnJS8ziJqk
4gx+zoCpNRrLFmUrTAM+c+8Vdzvl8yoDVr4hrjzPtDw3m+5v7Zy5ZOs0jkdo+DjL
42BY/eG/UNxhMMrlOflItwYwABGCylRlWKCVdB0HARb70/hOfRt9rDhAhQFV4uqj
96TUJDT9p6Tbo+/8UmUlZy+cmG3LL9d6RM1lQmZ1X39zPO4f1EMRrqL3ZCSZVcYY
e3AWHMX7EBefoi6fna33mXuOY0zurS7kHpT+Xhyy1nqAydjYDKbKOsfNYXJO1l1c
SCkhzofwzdxeYK+Kiu8iB+PCQb1+XmGkGBMNmUEyjq/yyD1yWdqB0AWOC0tXqwac
divAJpQWKokBhusPBlYh21EMo3mAIRKe+sB6UPi9iY6Gejefy+Vj4vRfb70Tu5tA
R6qR29yEADNhFXW1EWLCoyTiaMjnHWHcNG0iT7kvIzs/FdCPmU3/Ic+NvkF+W+jd
9IxM/rmIKnHVKSAD3iGHhik8HWJpabFtyn5nial3aszjLT/BpXWE4uiRkxU9IRPD
WdEWeF5cJ1Kk32SR2EvzH0ziHwZZk1+UWHUjW9D9racwOQgcNQJy19jtIBBOAaZj
jwqR5OgvKW4kU9wk4iKz7LAr/xqKmkkujoW4jxhpO0WNLxlnkdivzf/C7Y4VlC/e
y0xg+e4gVP61/3xLhaxexpjrHdc+kZsuiqjxCeCMDYPH+0LQ8/0CeggniA7oL3Ay
3OirIazvSGLqIOzNXAbdIxPMX+YJ5RP+QO9cYrKpe2+BKTbNZGzA7EHTbVhCEppd
Lihwv/MVVMmXDnWNHO5dJFd6vi8wwIU1FzdnQK5E/urFYYbxZxduf1cBkYZiA0+4
rTkAnz2U0Uwh11WaXVAkpkgCmQLIaa/FqUU9pmlqdprcR4s7bsFp453j5qN0K4Yq
/vRfCDizXvAa7B8NTMx4+k5MIZd2mtRkjWdz6MhEbgTGH76MasaTfD5pIMPb7PWD
JLeV0PPxnqPC11VkmwzQ391VS5jM/vT+9i2VkS5GvweWbPRb+GnbaVtkIo+CUtS3
eE2pzG6h5wPZmOROOPqX6S4Bch/3L4IxoDrbEer882wLROJy9UpZChpEldl0G5W2
TkyS+qQL1QNPDYwhPCPDPaf81GT5XFSe4oYqlW03TkOXruAc4aLUUFCXPuHOCgNa
WIeYwmu/PCbEzOkstqYtqNC3JwUU+et8Z0P5/aOOR4i0HkEAhlCXOe87VTGicKZ1
RVMmILgFT4VbkNoBEd1KL1iueKR8aWMQGhRh1cue/jwNyHtazkQK+s/dIQpOt8Y6
GL7CZET/Dsd54XrhBvE26BctwTU5BAR2f1GR1lqKIslCtMA4qnky5xY3Y5TrYUbI
gAqiuNpy6s3Yk1vJFOwaVnAh6eEVcWBYgzxtD04W8N2jjcGdXFmMqgCVWCLdKrJ2
8HAivOLvhw3IuzLG8GUvLnjzAt1vkI4b38P03Bb9vCXTUPr3wCtr6cXfB2c5opAn
e/ODKd2+VnaeLMZFTt7pSnfFVersmM1Z51Dz6jIb88zy0QvzFHpbPKGTCG+8FxdI
Ro7g6cgqT48Z2klNPoFmhN1BOTDLAWbrYOggn7ezWuSMGmIPxUG4PDwOQOQYQxze
17+pxPGMdI+QjC4hyL5Jbj8xbCJdN5kSXhdQosNrFWlNwgRnfZ29thvwMiMegnlg
xy4ds0gnJ2V0xMItMNDupMhjV6Hgt8PFmGoV27+N52zrwH+T/49J6CgF+5qpoiRI
XZ2gFayywwugDtsyTDHzsA==
`pragma protect end_protected
