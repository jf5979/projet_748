// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
0TWr+AQHE5fRVeVUV7vXH/f15HyVrPuUqryuMf3Cj6EPlHuJU7SAFOxVPesc/+ALkxkID0OlwJoY
8qMx6818DZcFSg91llJsd+2Qy+ms1SckXMS2c1wE1SiHdmwSGQBvDGgQ19WkouOOsfbpWPIUBFC7
9lNLXcXDOiM4EUerT+30yv4o3t5nJRNcCYHbu0oGkmPAig4MO15CzIg6Ivc36GoB5qA0swabbnak
TFvzcbJz4jvxFMZEXxxyyyUjUINj7u+DYbR+JuQ9wbTnmHJuHP62XJ1PbgotewpXZcuJ7V5XcVGr
iDCFY1pFGwTnP6yGyRWgAwJX3DpZ64l7twBezg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11376)
uBPfeFlw+F4AcGgWMNFnZGHphdTyNO215trJZhYuKkIn/5DLhuOyOckwb70Cl94tOybMa7tGs21S
p2OlCq0JS8evBdUeG0AhgHEdbLegb5TaMw7nMWuXTvdQIy5rh9dZOsN5Z9EGg2dDzFnll7kgyfeR
br3JP/x+msbMNho8iEB50yWRUSDpqIWNe+w5MLKuUpSya0DUXelW2Crc5AukYJ2gcuIYfkqi1W1d
vcYiFAbf10kZOmsSTbt8FcSXGbUgNj2d+GsOy99X29rFR8iXTTDHrZO8B0Xg0DFj6Nmm9qEKH10Y
+1R4j0A4nRg0wnfYrxETF02phHuRgQ4DNAcwRLSzpUJwhHZuR/sqmr0BZhs3fnLW4kMi53BxBks/
Gi9rhxUwebKWfyfH2bd+ykxxYYVhN3VM7NViFUjKfykbsZfdMtLz8gmxpQEVi9ZA12O1yN7SnEM0
UoYf4l60/dVbEPtIQntJxw3Mbpg17vzegyoCTnpUb0KEJvbhKosEOOEmm/2ZXzzKGv9GqXg1yF0p
WnUGa3I+p4ipsrqwj+16nRLmZss9kCXl3rq4fdTZk7p3Xuv/T56ye1csj1Z1ktDD0KF7zKHsqC2j
/IA56Z3xzfqYkSjA9sRKMQTAduoqS/yXv7LO9the2RKJXsTNlkc9zLqpZx6OWvA7dFQ7rZOCy9p6
SNZXObkivhXeRMCd8uISgZqlDYVGtidjMyUcbDbTKpuHfa6Z6zvqFwXJ1dueCAWiDtow9k1o70MC
vkFhUPH9itTiroeYC+Jj9yLLNlGP3AbsJ7YzrnnuUGE0HoSHopu9Z8SQUMfvGJOPu8oW6pF446n1
oY3sNMx5w4zwKGmU36F3FxIIVxZgZ5pRxO6eDSGgkQAWvuRWk1Supex/hrik8ivCwksNpxyqUy1f
DSdaD1fcTKDotHKrboZH2hYAbXtpuH6C4/SFwRyBGhK7AsL4bnOL9oafjeZrQhMKLtyLldy0lySR
TEcpkACpCEnia4tl/Ugbr+WAA00lwaJ2GqtohYOixKlE2886FpiT1nsW11A7SBO1oEs2GdHvQUVO
iCfnTeZs7NcKROJwhAP6yT6YNyo2cdM6KCsDq8nS2SnNveE6L9X6DkGJaxTNK7kq19MnjF8to21F
0Of2PvFO2xclk0BxracRzDdLDJX+VURaMMkcTPDRHgbOhzcxobRqr0g5GZWyAA7jG4trTrkI3dWZ
HTVKljHflnLKbdvsTa3oXiqPyY0anE8ORV0HBzHZKFdcJGJRlfxR++F3JujlDRqKjAaIiksybBjd
+FwDaBxqPZnBNuhj3XsF8YM6UGCt0cmjXLSS5bRszmfzeDkGA2ms5mT5IldVmcD74Fpy7GskjQG7
IqAqAgN6ifo2CSeDr3A2bO1Jkva3d+ju4VdwxynhTZCZWyHzA7n5OKOW1e/AVbHU+HL1GnK1gnxJ
T/DAd+AIpJWeJQlhJPOkAX6+w/kl/yGPRRWkD4XC4VdBzeL9DmOid26rxVp7vhisy9uyT8n85ZXh
564RV4rchwSHL/00nGtBEqkUCM3dQby3+g2nMWjCw9sabMsVYKrQM/Ms310cWHZtUZMe2kTrB/GD
4ZqCPTbH5RrwFb94sSl0sEA5YqdlxbVA0VyVRajsPMSYmgOI+vEqlRgiW11SlAlbAcWQvCTsttFH
Bvu0FMY+KF9m/Tsx85PIyg/d3/hZeLvIr3uW8FaOUAOSzsKtdOw4QIJ3VrhLkWXOg/7mPhnrjb4e
KFPhT2uXzP24w68q6NLV1VskwyCklZQOgSNMVjRStjhiAzUdCVBTID7EqgyUmeS60dMpzQdlmE20
85CA8X+E2aStub1luJP3BaXh17ChH9tZ4rwxZNWcP6gAMOsJuCUMdfk/loT9fT6QSaQMB3zJFrNP
rc9C9fOWMDuTeQc1oNLqzOdzuYxO0NSSA74iVANJlUmipvChIlnnekkIS+jM23G9P5nsrSTKOEf4
edUpeqn4t91izIr5oPOAlZBJorVHC9VHrTwihbXSBQC67jVwf9PvPBCtq627d2dfcWQRKjHTaFEL
+JqWK+HqAMvVmVxcCZKmSE10t12e3OiamXOMZFFelzrn9TwfBMI/l7mNjXT4Fj7ymORWa0rZePmQ
HvrU5U7P/6Ez832OYBAe6wg96ffjCBLfts5sCXRyW4hJP0iGXfEz5Hpw49jbbNJ67fMcKl5u06+i
fFANVhK3hYYJmjYPcAhNWc6v56PClfbchyiV9f4SpdPjl20e1J9UwZHaqKBoT7tOzTnSIVVZXDBD
n9DRU/ZeiHPlJz6yNBvuzDoqjPL49DBrNtdFsNNO1XCkPb9sEl8znvG2EMF54z0W+AqcnDHTA6kR
3O+pmSZT57jlR3hzpf/zEvzHst92Yjahu/sI+id4B2ykn7mNYvzvARyx5jTozeRNE2wHNUnJTdlX
lmqotkEsU8+ja+PNgpdEAhs46xh/JsRycfanqHLcg62CBhKzoMAUVRzbcrjjI4+JUtnM3CcNCc26
t3XME3P2ue1Lpcb1D4Hy/Myn6nwFE/0nUGrfN998meUxoYe33caUBYjCk3P8f2BHwiiuPyTKwufK
ywxmmBVhCMRJZhxKJ5+P4mSji3WPlZiQk3F3ghErkCNFsSO2jwNo8KfSsD77PvumzaPahkUFPZ6p
YgOCvRvqejbeYsNGig9b7VWpMVJDVzWgRpZBytKIMCY+KnQPBvRnpgmRabI9W5PaAM4LaV4YcUnv
tfTAXGgXq4KDGpqDt2NLaOPzBWLDrTAQcnc2Ja7RZ0B+QEFtywZKzOhifjkHAGzqFzoPgXe/7VMf
A1mVLWImRzutNKWK7a5/8BsuK+t4ifoK4r3tqpNSU+CkaXsSu0z2Z31EcwE/nD6HrjITolXiI6Kw
7lz+axNzt2KgZZ4snxQnEYTKdx4ingbehEInPR+X+v87Tg6749VsL99D6A6XSfpV/vziwCtDTq6/
bz77ChccBPQndXIyYhPoe3LArZ8bMyWRJbEzQhxueiE3EkSOMC0CXGLCPaG6AHI4aES2dbQ0rqH+
0A3Rg0RqzvcC8BUUD6Txm+QxbMLj6edrXYZA7jNy5gtJfmeGU2PIhtnqpMP1O09N9oEYpDRmBA+e
J/WEldeF+7QtMGk4BtU3euvev6MVM7LjeolQELOnA3JZrrmLIALVm5d/wvCxwLkLf/knmN97ULIx
XZ7Rh+1FLbOtcjPUeBXeT1+molK3HxqZOXCtAglFE89HLqB72j8Oe444+8EgAJy84CZLnFfzr3m9
xXAXN3+N29gOipBtpUnAeMAJhvblzwFidbgZm+G4p8pIYplun/U3DNvhuBNBVFN2DyUp45MHhXze
q1QA8ODYm3fo//Jh1qCblJ+lHWfyR5QFQf4IWJCunHLyGMQM/K35D7Xb5mfLgnu+yGep6OYI6eKe
i5PmVZpHdc/D54Fj+0TtWDrFpqRFRgsHMs2ZvToBiwlj9gPI/kUgXo+nWZBBs55y/xbzP8ZRv5Zo
CDHzIstet8GWjyoReURRMvfklOAlgtGlk07yNH30BOIwySu1CW9HTv974uevksWl7IKNj/ytaQhG
EX6ouw2/RXmq3KDEJE6+K5hHjn2fqlGj2DI33+OhAESy5YEmWhkDQFPqc91mUx6f/bjrO/ypJkX9
Jxxu8ZLZTn09ZvTHasDYKeBR8W4Zt4Q/nTMwGfedjaRYUFJiJKTzzMpawefBHr2xXK6G34N/OTx3
q7RRa7Uq9o8E2KkUbwiTBzRjBlEZi1/rt5VSxQoK8jZjKW5zDmjeWO3FUagY0PXHqmVZvCpJHCaS
LJjUbPtj6KO0OZYWjgBbU8D2JYrwNiXUg83PgaJsdEUNf2mKe3Qh5a+LpaFJqXpgynq/Upzl3WHa
QgkUcVyBEAflwYVx1OlClaOP/xjfOLJLI9yYBkja2Nbum6aGmggZl7/z4we1B54bmSBkvyhdairS
W5VZnn2mA2Mc8n0IYYYdsuSYN4IaWcMu3kCNNszwgYBrEapb3RQb/4e1Q8RyvGvpvI5qlxCPkwmy
+kjk5m0J7GewOnebULPJkS4tq4ZTiIH4lfz64EqU454FFcwshi0VrMkq2opCOVahcO4DdjyV3yFb
7nW6nWcM3hr/1eEqCxtLmqPsqfrwN0GMiUJKy75S9CDg6Gvxri6M64HO+AgyMQTJiZLHa+8Da97D
c6DUZiTfn1ACOCve/vM/MEOiKXoQw9MZs6I2n1jxBN61KkpSHPZ5Sb5lS9rljyNwiIMsBW/Q6+0l
SzCvPzEWGeR2+HqdjWlBA5YgKvA+C3Wm2GYUVy5MAh4T4+KugZw7JH2ZgIrzp4n0upg6jMewoKPL
YlB29G2jUcWMpebfXaRZ4IsmInKZi9Pgz+gU8mQ3GPvOXuGkIuqaugo03f1BPUNWnqxah8TJQjAk
wSoWs5M/11Nnl66JGHr9uL13/QE79PnX5fsxsG+qW27l8lfI2sv2Q1u+PEPhYvo/PuHt3B6NOS03
fLzutiUjFyfD+ZNE17JQR98Rd0GJv8Kb3Qyyo8WralKWOFKazgHqoZZMVmGpsuI/AG96kYggkVwU
wqvfXZeHBXtkax1KY0xz6pY1g8lH3N10ow/j3tCt7iUoftVMK2MOD1GWzy5psxEqarmSMV2VrxWg
u2GEhk2iVArpKbvEgKPZxaedmOKvqnkTQimbr5Jv+cKiAOt+3pt+ezQJbBsPp7eg0z5gNXNfpZiU
IkCRw6lj5VYmDjXVJMT8RfwLYvsk+Zptevt34r2a5pnlBNqbaNkHB4vi3/uqMyNaz/QRblswhKGc
smfm8StiGZ7xBAe2n/ZMWFSEPNnoqZPDpfoVi6oOU0fvcN76Kf5XwP9fUuu0WYvVqliI3H/8Fq0P
SC5erYhs9Rws7fFvWqvtqdoqaF+ko3CpHIEDS1hB9YGQpXMKNR5j5u1w7+bNvSZs0bME13/t3vEv
OFQj3CGDhI4SKby4kO8rGGQqcx61R3CtBokbVZApjhfADPX7kTRQYFwT4GPusplgQU05eWyjS1HA
OOL7YfwASKyuG4u+qCRQfRDVSkNBrOfnMahe8diUfHoDFDTSI1gqsuGB+eMhxDuy0qx2tA485qUG
J+WE9jkafsMby5NjlLVFJuvI4kGydeflCe/Qz6jYSm6+dzYwRaaVEimjc0h/QNluYZ/A64tZxtTy
NJaxzpmVnFOU9Zb4+SK8ggihCl9FyCf52OThT6tgIWtYnToIlPqKzns3RvHz89nbzq7RrEZ9YLSv
OIlhfbSZL3O9nPdk79peqGyRfR/CNUEZoi8ixmOefsBpQs4iEaXDquoOQ1xIlClx2QE/+fLIc9gX
wyHgwlx2m7ksaG74u2PIUAyjs+IXmZPgE7js0/gSRC55dyV5RjdbOYb4LIsWyS5M8vwwQeCX5yLc
ikxrmL0DcHXzuTe7eLqncf8m9kmwCE9ZJJhvQXPI9/9Kvl44vC08FooX1fkYZM5sWpBkEe6TVyK+
0HH2xyW7zDJDt7y0CE8ilSUP5VVYjfajBE/hSkKyNn1SIvcdo6WY1YGlTs8a3W0aOeDQuhZGubts
v5pbRGR3D2WW8VUdt1Ui4nWybZV7OkI4KBA68XQxZ+KWCp0np0PnPVYkxrCndsP26LjV556CxP6Y
k2JK/B45XB7XZq1lwdx2X2jGmDFEWfnRmuMpSd6Meqf+UsBUfwpmyvfcOSkiItf2mtOj2tXdlVNT
S8QvK/Cdz4uJRaZ3aPspanOZDrDv06VIsV/p/HyrC6lc3aADk9s3fNITbDE8p9Pm3nScUqeFPHcl
jd12qANwovtgzVjPiJ3jr7MF1IyHrBAZMXhf4Sukr3qqTzVOSCkypDNhEkFHJE7emfLSbjOODBRa
Zc+u7uP5GpMV2QFk1ILoITo2BjtL87Djo/YwNk87/jkA9+6Z9Xf5ErcORcAjAHtygFZL/mqmjHaI
6VdWFrgAe1o2YZvogduLBtDWw5mcA73qM0RhLSXQOvOcJbrHMZMdPZdSkaPyRTPO4xhc3XKUzO4M
PyZ2zNUi5bebCiuecJgks/V/z+Ksa2VFZ6mJVYTLhwOdvf0PyLx5Oa/CcqDvUxr2vPeco45uW/rR
AoPf6MMXrKUf3riVQKDlWBfvcl1LtuufwlSaBu6+R3RKeGxM+t5i7RMqoEc8V5mCrjHzNnXnOI2B
LV6+Y2z62oJCHgl++6kOsf5E67Cr6FKDNxPv765iyySqjUsRQDF5OZDBlxteLkQOy02fP+/f6+lv
IzjhPNFKAIhrBgxqn5JqZ7/8Qtn0a1ikHx6G4PN63FCTIseqW0R3AJmDpktkb/wZ0cuvQT+TuDA7
688J3kg6reFJ8k6KfWhWGNKXhZw+dWckZR5e6T3LO20ysWkpXCZ1ds1DiWyNOfCaOUUpaxzygif0
TtmSrCugYDzF6EucE6TAavMjynEj7BREOGwMbzIRKDd3qpwVgZeeLRpFGhrmK3p5BaCy1POCBquG
om7pH3rZhe5UIqyUtXYkkHgVgPaCrxvhXCkCJgqGTds8Dub9OwAPw+kPCX06/hCa/fQMD0SVHgSA
6nCZ2aD3Qlosv0rzRo8xxOlG2JHTja8aF6s6cE/dpYusA9/tCHm54uGOKgpMAXtq0dVbQsaYgigr
Dj7hqS3bEHSZcldhYk8pwGnem7aJrIel+YxMQGhc7o7kxvH+difJ6id8iMHhtCOdkyag4CZR/DNw
32sWa9XmbXf+Ft1dokjgVMKrv2IxsVl8slBfbzF9C/azX2EydFpAjtrzP3fAhlJKzRsbXNeevCkc
WzntVo3w3zd5KphLnJvxgvWDdY6rkJPCxqR2W65gn8gJnPW22Y14+uD34K2dHmHVbg+7MAHzB2eS
CIkcXs3dJoCK/ggubwgaaV+fhPi4+obNLxVIauHw/IhaQJo9AJXcGwGE/R7WUxHoRLY5aH+1nyjB
JM3DDztxxtxnJm3zsfyVVLgoHGP1M0j6aaW7rZuL5mcU2xjdgTmihmbFXxG8KdHsz9+a6qh3AGFl
+TL9OY0lNDFrEvXMa3zTdiHHYQkgrRU0fyT5u2RJSz8wZEWLoP3VsEOKteVy8xXnaAhNLdrDauQt
bOs6k2CPfOWDY+yGlvw3JxLyUus2hiZNA6Hix4C0yHcw2ML7o4BgkWwWsBIgyKvgoYAlKldmKHW3
q71Anei0TAYxRr87vEeBFp2tN8NzJ6Lzd+z16rvAts41HPw//vfs0dR6ljNI6NyVNQDAJmo271fy
wUAxGarReDmpckqjm0s838UG14WBlnjwwtFFor2jDjrGPNisrd7WhXBAgKs4fFUmeQHqtfdDdMUN
p4ncneasQg8c5zQM3x8TVGPwsWZtmePrhU8POMFlRKML/1jsegTbQ8QWf8N3bM6FovMGoUjTHal0
DFERoCDu0vKTBOULVnoJByrOKYNfttJfLKdPaav8mr7LPbswQJc3Ttzkm45FQP0jOKIgkF0g/S9R
e0KzxnJmp871Hrf3ARc5wMdb3rBOhpm4kuD1EZ3sL0tl6YeE0DqbXmVOJpnl8IUW6W9OW9dHhMWV
Bad8qQ5Dk9AdOj7iW6MX7IU3jFibGRzw9akrlsi1P6UAYuVabgaasS7gzZHfsf7+Wm0zQZ6mfaVb
y3jD+A8G5DzqwmsXwi2q10MoRya5fUO6YPNhq8eQ7PDUS18XdHaAcTdcfF81P/ZoPEZrJIpStekd
NUgSPmsLzHnaknG0VQBJDedzxJbqRBjZ23/zPvcFGlFbbrE8DTnICJOHnw+Jg54TmgGvCIoMqkcn
kBV0VDVCUy94V4NwI6rBYDmbrdAH5ryrYU7z9BE5mq+GjxHGjQtdx2FEwh4AHOzHDIEZQ6+dpo/a
V2Wa94AVcBjBeIoywQl/KYd+jbJZBCc/rfGgESyMGKtujvL90/Q4VMs5mVg0ahGKQ6bYD+0UoUUe
kh8J/e0uPJKoGzAOnyi6/UDZuUjQXI2Jsujp/U+1DuUUiXgdHxtjv7XAmTJyUfl3igs5O8qPrleh
bghyYWT8nnx4MxAbzzmqEwgYqpS/+7jBokLVxVL0xVsfIN3c4bt20SNJpxDpyoZ94JNWXu/fFeA6
tIlantb1L6CtK45CvywzLUOQssxNSxIoRDOlov1DsKcnbqj5z0FkJURNGZ1sbh9DWxoq3KAzmzhx
hQEdM5fX1zmJ3WOxOe/edbK2cIGGpkxoojSeLTziY+EGDhnnSYcJLe4whY/+AatWRI3nTIZP1kHz
00XimyRMYbIquitb+dgNTIvnpXA7dPTGBkG7TiGdbMavnzrlrkItf8agM7VTSt2NPZw0Ti9M1ePk
40EBaFO/k4jP2tZ8+ENeCMMboFTVaX4tnA3iK7D3m9pou0s5kYjkqeeeT//ozkYLwj9OK+IeL+Gx
qie9FWLMEa/JERr7UGCMUf2SdL0QqXNjeyewP//TUjpVylU+rWLgYNCuYww7NmCYQbQOfGOpg96E
Q39w9C+olunox4Ab9u75MkMD+EPQjNZKib1etHqWxul66avQH5BqSnwPJSY3z/OiwVEfMi+lbFa0
uUNdDgNsulTPJKuzZFWG6x3k4uwqIJxA0SO48T9HJNHI1atEcPhi1cHxzd0htMgga80KgwNde/k5
/ognSyZTYtJX2H2dE4iq0F5XXZosOoBhIMfzcFe6rtntq7LV7G3AAOhF3zlKHf5riwc3kbj2EEf9
0pCu4xI+NMuheFIrkkt42ylof28n93Jl1wXvORscLC7X/riMOJb0ukhzeySDWxdkuIl1vrWN5HZx
Z2au2/E4aOgqV2HEEnCbSzorRFiGOf68AH6mKtNqkymnaKFsXwyXYlMUJPbCc2W8xSbJRWsp7WEK
JlzSeatJUrAJET5l0vNxTRK1BeJTSk9a4J9CkkPipazCuDYskm5vCWEIlGtmSgH+huDqrE6slJfF
vIAZDB0dK5lYBBMeL8IN84Ye1hHyqZ5/VG8luOW6QFJzREAWpg168yS0/ddu41hGP6nSaSEol8vo
6VYvTY/iBOio3UcgSVV6FKZF8/3OnFpF1Zowy/Ql93bwiTseMbdE74dsKemsjz2SiY7E8DfRp2Z2
QrAs95Plq1owKdOL/ujEcPCvvryg8h+d3tQEqdcpn70qvrlDlIujJ3xT0ZcAhIjG6disAj/OJF1f
fRxYcSnjcpCxp5muc5l65Hm9o8sYQ/0egDUacEtyQy5avi/InSOlloaKGiBiyMYS3FOIg7/K6Wao
qdcQno3mavEg4kUO9u46BUAwXutvQw3X/crMG1GKnuKXnYqVfx7ko+pjGAKcqje3Yh7Z4oCYLnXg
QNgGdDnCNqKTYaTbXefO3wpH7HAHpddhwk43r6i5ZTGMC4rR6KYyitsX8RwUOGebcXGsEu0TF2Te
2Nn/saF/7yXoMrTMcXQO9wAs5ZoGtMxDoU7wr7zo52FNbI2guVtdojr4wMq/wnXTSnVYerwIEIve
HahzZ1GlQ3o2TP109uOvIx0+jj54Ytxs995g4cJHxMmsD2Taf/HHlNe5cj5gpq/ICOZWBb+Ytn6V
v5JFyNni63qvaKRv18KqX6CabwBqc8wHVuLa93/XjHXfW4HNpitRWssM/DFhLaXJBIClANUhp+wU
m1uzb9wRWoBDa6wxu5gOdEPnWOhAWdUUxGMA1JaSg/jsFdhCz9tN6dMkExT0kH5U0K3JMiIbAkeL
nbF2GFQINh8DuyFnLb7+tQAtrh6DdxaFLXf4ekfrXKkbFO+QMyZ+l4qKmrdbRAZyNBKfJB/2jOgV
Sfv1NqcP2PYXAGmafnE55RqunVq3wWsqqXgh2Uqd/mr8NUjCnK/0IN1iXN9XPXIUPrm3xgMXn+fj
2eGylVA4PoiCni40NNC9r74naq12/u+bblH2NVV6E5qnfVYsCAUwWsU6+KOV+U8BOeA90akH26rQ
2eYHZnCTZJ8R2jGCDc+fy41C7wOK0mLT9lbM8A/ZWkhNxk6ZQ5Lyz/KKfbMga1O7p4yJeuJ8NIFo
synWUGufXZK+d+CJrEMKTHs45YSYNy5vRSafW2u0cNIpR+eKDt4DIVAlIC/3bVPpzZqatdgQYeVx
xPgvSiioex0vPFQgg87pJHO1nKV6Ioks4IUoFoQBLTsb26oPeYT1fnM+L09l5UAQ8kX5Jp7Caxkg
D7mhPuOTl6mVi4900lFrUp8lWnKwLDqBUEoRWlgZIOvId+4BrZSqTFVpj6qEHKu9QNIphHJI/3si
Sgu8xuU4wgZ1UDsxKHf5/7Vm8jIWZCVsMOL40fQlzd5BkwAHeClM4nfT2MaDI2wUyLEioixT3OdT
i1+kCRz5Jwp20Ht44z4ejeGzcGlQlaSeI89PokDjhbpynRPBiGCPPYZ58UjGM1ULVYY0chPj/qX1
NHbXgD+6z7jgSu9+ofRXmqOoBSmbWaNG/lc8LkjyP7NaCrHLV59owy75n5t9Pr5bPyEUJ45xToBJ
JkcnPyL3odQoGv9J4PjwZfpiIWAN75rCn0HftJeTdMQYN5Ah63laHZEZwEPFdahPCvN1NjNcbGzr
bkBp1N7ldDnbdC7ln2kvXdZ5gbpvH0op9YsW/YUtiCCsTFwZFeqTfG0YeJjz7iNLM9Ui9c9t7J2v
Wg1O244QkncBHjx9Ca0uf3+LK4ZH31ojH4PU+Qjl4LJkD9/wHKMXsheRUlVf7euLNhW/26WAQjoJ
n7Ki+N0tNaTMzVUJSyAV7FCdaK55Ar3F1BEmIZqiwhW4GzyzmzaSH91OA6CJloCzMCAeefMoWsA0
3A4UoJhWTi9W9EDYEwHNaVd01rg+NiggnNNkr8Ac8YJd4IulMIVYH7MUNuJT81/WGkmqbDmXJYPG
N7hxsTx8Q59fDwY0AgYCcYaXRoVhyF1lPZlLxdnrBuHcBKL93wNH64Yg8zTn5KFTU4bSJmIcFrpi
Zw40KXGapa3sS8mwT8FmkwnzwldZV0QkvVewB+nBIjgqSh5hY2ZbRdEebb0M9yUlWZ7emO2poZhI
4gevyair5WxvHdk4nvi8gJM5NIV1455+dgm4KaWeOzkAa9QrfLhzDOVeJlTfcoHoLucYNKyyySP1
RyB2HLOWUJFGpfIPlJmWtuU+BHrhPbDFFlNrs0PVmwo1h+oYqzdcVQLOVHOwofW2KlZUZ/FLqefW
ei5N9r6I6RPYTOcH7vm0waLmBOSEcO8vlTKzpgEeLxlPp1ZhK3RM9iWdZxOUAqYtOsIRBh6IFTqc
AI+GvLTK8Rj0cmz8XTzJ4Zm6Q5JZMxv3TFXeP87GA9ZcNobJ5U9/JOJSE7Ti1GnS1+8N79sWq0jA
yygc1Mkk0LR93RzoNuUjoDRb6EHT57gFfJQi4U1s+qbCE8qFDNYqf+jY/UUIfl8b9IChznzFUoA5
J4M7Caag4WmJ6AsgaDE593fSPmIJXWETFQRAImcaFmwTnBhkVk6wKwq3RAroj2KCO4v/WK1eemzm
HLO/Ko5sgKHA0sCyJ8b3sQIIlkvAlMymqG2qTqhxZLBU8AuhvAkW0RHruambRj7rw2480mMEeUB9
lDj0etHHIlIpijip8bRcTalHf/cD2aUhfdz8ayVoA6ZDx7+ma4LQXw0F9dhl5YeDadu1ofd/9DuY
X5J5tkwSoG6E2W5izb7boLGc1K4/NgvKlYLWCtU4/5GkL1kB1XFn0YM6Oe2xP5Sp8vL0NrWJZ2BV
1zO7ijEKJK9ap9ubPecFFHRS/8WCwhY/WEXvKe7UpTfCjpll2Q6ZjJR6rfjkpkuXyLqrQmMxuD63
0LGVy9+Hz56F+yfOzdoXHG49E6tm4Pl7DdB38U8ol5D84/fV/rBRMIoODDpbrxoe/tgEX8I52YuJ
i0f3lMp7KEdJ/GZ9qq9fVhL5RjOnAUbWPR/4PjL/5syeK7WJIuGyM6PnE5b3REmJXLpBwBg5meiG
R9JCQ8gz7Z/cGMkOc3VW1OTEeDaYlIN2Bmc7zTc3svW4SXm1MJ7Z5AjDlX6EOP/7CbzJCkzMBtgS
L3YcQApjF1au9eBk3iw98ElShjivV9FmgOJbP7gJELNC+IjncdQWYr+Edybzs6lP5L+jJ898TnGS
9RwMOvjkpH1CsH8o5585P1Id8CId7MGenBNXltMWgNEDL2T+8YUZtg2jFr8Doeq+8YaSCByNe1pu
iuoUkfQ9f/+uLHId9cjT8hf43/UFN8BwmPjr0QkzIdipCCjRmD7YEBI3NO/3+PftNVrVLYRUq/r2
pSwJCEVIUKt6KDBweaZvMD64M/X1qFkTxgYyAxYa5tlv9iiMRh+wnLewr/oYzFpfqiXZm973+yXh
P4BU22zNcznlGQtaZfwDMMtDcVihq88OioQOufNMYg1FYRUHQ5fHIMASbOJR1RDPgJNI11/wl7An
8+lVd6pbHhc7nFnFqzD95re/A1u3CwaN46EYqteWJ5qrmAx/vjmGf8wx2UDiHj09b3eukQ1Bg7KW
zNfImHA3lwLKuqbWVa3fxh8Vp6OQ3cM3LnKzhuGFs9+tMUk0q+fMZErb7ge3B3Zq13FQ4/Yo3VbO
yZW0KuH4vUC89+djjWUYKNV2wGGTwh1Qo51VYOgOiCSM7ieZFwpk2TEV69xJYcpxkJBurc2TIIWM
yn7qSWP8LK/leqYtGL1eLxFVLJU4Y9NkAn24Y5gUEvk3bU/xyhOzzmdzOIK8YRX0UeWQpTEVu/J2
JZh6QC4778LoqJit2QPT4we57L3iC6ahuFsZtuMM1Uh31rXqqpmgR+fDngRuASXY54ALZ3jLKkXL
5bznuiyiQrJ2/ayXZemdMtEaI52La2OGkT8rJ0qZrswxJOWGdIPu1arBnkUAapHk/1R6XM/J9iO5
YzujEzTeBnGyXW/+CnzMcFmltW6NlC4+VIS58XEaG1+Q0Li3uOmJT/Pbtp9nssryQ08avklQgBMs
jv+CatTi9sDqEHw73VRZ24J6Frll3F1PQ4TYjOHTq/IuvssZ8EU/rOUWUX+agD7e1qCj12Q0cdwK
niCbwGIgdm9IxrR0ahxeM/r3RtLgCA6QasPHUg/l0CMFocWwvR8kw14ljNyItYV0U3OdrCJb9nxC
tUfGqRHBe5VT5A2TUOGx7+eCBGVu8BsGSFMAfLS9ObmkM6BxMg9FIzufGyK9EMp0wUvgaWGkbBy7
WmnppRYgplRAFhzGkNEYtNaittkA2l5EOLQxTQNGnlIJY2QV6hCtUSkYi8SckhSCw4xRMkfV2IEA
PvT5mCINZWfarElgXvU9VZAKdARyt4d1p8PHFn+ed7DKEm06W6uQafHqSPzDFLGMraDpQOsiv3Hu
wrKyMvOYwN7yiQ2UfuXPhOepsv0riMOv+2AvAZxtkL4ww5kcWYmLiTjuttcifMarJ/jxKkBt5iGb
YFxQcXoQHIYHbF9ogyvzlrv2n8mhfCY0LrXyBI7aFlXH1TurgzEz+E3ZGn+GlKy9muOqM8Rs5d4A
WlmJjQyQ3pR47EE9lWG1XGBShIHp5Q272EAB860sIbk5cNwhJIuIS1lXO+A+oI5+wNVDmfhlqP6T
BJuwNFiTPEkWmp69WXARZ0InX7RlVT7n/s2WXVb2fRNT6LAeT9YFTUunDIUMjNbg/r6zutrYfCVm
OwxE0FMW2++cxM2DI8qBErLOVkL9aZ8B+NfUejZZx5JXaMziYsM8eYOxhpZlnY95eSq88pWGb9Hp
Mtg7xNlUzIDM1CaihxOMXzAOuC8wW2WoYu6lMzuhcOAZEtK1dr412PKdKbLQ2nMp9cWe6FEvF44v
TejzJaaNUAnrH7TTcv8OqDYBKPUvnEiWms/cQYOixz/QjLihdbpALquOI4vneFsuLJ+WJLj+gbL1
VRNx+CI6IRYT+kYejsmAIz0nkfZhRKISwb6qVB1dY7FDh0OqtY4jKw5cl6t2QZ4en4DpdnhdrRQX
UHcdxRyL6KPCqDPYsQIhMkcFE5Cl2/Psruirif1/RWO0k+UraPCuJukd4BYd/U8KLqIqEH9Txa1T
nC5iqgRVdYUCVDm+dERcEWvWa2nnLSR7HZ5JhuqFDX4lrv1XcJLHHkIx7x7z9hmZbRXwwbUDccT+
WdGxaOj5K/e68bZ2N7aY7/7/mS/s4VHplsUL0IL76zhy4XUoJbNKnBx8fYKUL6AUwjAkAFBy6sAa
jeA5TsWZn0xA2WgWXBoW0NMSin6VqDK6vhwLk5rBFpA/LzCBjF/Dre4LqoVgoeUwSJ5I0sKjKVm8
NT1vIODfl3OxKQPGBHSMWprKjzDn9c96S/vBAByMPY0yFQF809/GXpiAxWHeye7aqQQdxPf5OIq3
z7IUreXQjK7NMxpROaB2q+d6PF8TBheJssdiJ5/K9zQoloyIGQ3IgXr5K1utGR7RaW93eOigCgfC
J9U9ZemHN9nGgxacBpUhOZOAhsDzzNwOSbpP+G5Z5gJMVd0SDKJUJHwotfPnXWjzTMIGLRh7HFhd
0UqIzKta7JhzwmOJDvef9dc5hY5kBnrBH3IgGpN0n4IdzoOJPDZV7PUKr+v6i/V3ZxfvRYCnf00J
QrpCKVZL/SHjbe/GaQgQgCR1RBfgXmX/vTyf6ijXLj8FF0cRcEmd3DilXSndKpHa6zDfWIaSpkxL
QgrNjOHBN78nrmi6IJHroZoQymA+1dM9Px/qCzd/mzKV5Xrkw40npUEnzxoC2UVfdiXB2xPjfAt4
Zwv1lpCjHJGEZ6VFQqEbs/eEoyPPDL3VB3pWWvEONi2jDBky1KoagDPKdrRmddeQuNJ0mSKDmtwB
aBr/sEnqLaV7iBMuphIadMZ+11sULEVPL/Cbr7wyehX/FB+hHXCJE0Nv04ZIVSUh0nypDJ1KSBPr
0U2O4ugOQU3I+mjLvqvRz16h9f/vVJ+gM+bGyPMZloNOo46cIocDt66co+VoQgbEyNnfArl3hpOS
gXqLLLXRmujnb5MJ9KswUjwsm96/4MTirybA8J2Vkek6V+LWbB0s6Cgf+z25KFqDL4aQ+7onTcoV
Z7lEQlWK7bnDdQAO6qsYjybJ6tJb/yJgSUBeFMnZagKasEMY+iEsN496KbMmpz7HJ1GToIxLYW4r
lD4KcUaZZezd6xmyAHfYrgiTUHodJPkuL+I7HaBuUZJ+rIQ6TMKyhjtEaLSBBYyegrZ2+FmqDe1x
sPnDyFpZkIJbk1t6Z4zIPw6cqflWsUsWJ5FyTqK1vVA1CuO7YFijAsegJW2qktHeCrfvdmcM3jmv
mOaM27njiwa6FdOUxkv7sbHV74SouMGjKLZPjuy+TmAE
`pragma protect end_protected
