-- CodecAudio.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity CodecAudio is
	port (
		audio_i2c_o_SDAT          : inout std_logic                     := '0';             --           audio_i2c_o.SDAT
		audio_i2c_o_SCLK          : out   std_logic;                                        --                      .SCLK
		audio_o_BCLK              : in    std_logic                     := '0';             --               audio_o.BCLK
		audio_o_DACDAT            : out   std_logic;                                        --                      .DACDAT
		audio_o_DACLRCK           : in    std_logic                     := '0';             --                      .DACLRCK
		clk_clk                   : in    std_logic                     := '0';             --                   clk.clk
		dacchip_pll_audio_clk_clk : out   std_logic;                                        -- dacchip_pll_audio_clk.clk
		datafromaccmat_i_export   : in    std_logic_vector(23 downto 0) := (others => '0'); --      datafromaccmat_i.export
		datatoaccmat_o_export     : out   std_logic_vector(19 downto 0);                    --        datatoaccmat_o.export
		pll_0_locked_export       : out   std_logic;                                        --          pll_0_locked.export
		ps2_o_CLK                 : inout std_logic                     := '0';             --                 ps2_o.CLK
		ps2_o_DAT                 : inout std_logic                     := '0';             --                      .DAT
		reset_reset_n             : in    std_logic                     := '0';             --                 reset.reset_n
		toggleaccmat_i_export     : in    std_logic                     := '0'              --        toggleaccmat_i.export
	);
end entity CodecAudio;

architecture rtl of CodecAudio is
	component CodecAudio_DataFromAccMat is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(23 downto 0) := (others => 'X')  -- export
		);
	end component CodecAudio_DataFromAccMat;

	component CodecAudio_DataToAccMat is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(19 downto 0)                     -- export
		);
	end component CodecAudio_DataToAccMat;

	component CodecAudio_ToggleAccMat is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X'              -- export
		);
	end component CodecAudio_ToggleAccMat;

	component CodecAudio_audio is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			read        : in  std_logic                     := 'X';             -- read
			write       : in  std_logic                     := 'X';             -- write
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			irq         : out std_logic;                                        -- irq
			AUD_BCLK    : in  std_logic                     := 'X';             -- export
			AUD_DACDAT  : out std_logic;                                        -- export
			AUD_DACLRCK : in  std_logic                     := 'X'              -- export
		);
	end component CodecAudio_audio;

	component CodecAudio_audio_and_video_config is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component CodecAudio_audio_and_video_config;

	component CodecAudio_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(19 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(19 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component CodecAudio_cpu;

	component CodecAudio_dac_pll is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			audio_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component CodecAudio_dac_pll;

	component CodecAudio_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component CodecAudio_jtag_uart_0;

	component CodecAudio_onchipmem is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component CodecAudio_onchipmem;

	component CodecAudio_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component CodecAudio_pll_0;

	component CodecAudio_ps2 is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic                     := 'X';             -- address
			chipselect  : in    std_logic                     := 'X';             -- chipselect
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			irq         : out   std_logic;                                        -- irq
			PS2_CLK     : inout std_logic                     := 'X';             -- export
			PS2_DAT     : inout std_logic                     := 'X'              -- export
		);
	end component CodecAudio_ps2;

	component CodecAudio_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component CodecAudio_sysid;

	component CodecAudio_timer0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component CodecAudio_timer0;

	component CodecAudio_timer1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component CodecAudio_timer1;

	component CodecAudio_mm_interconnect_0 is
		port (
			dac_pll_audio_clk_clk                                     : in  std_logic                     := 'X';             -- clk
			pll_0_outclk0_clk                                         : in  std_logic                     := 'X';             -- clk
			audio_reset_reset_bridge_in_reset_reset                   : in  std_logic                     := 'X';             -- reset
			cpu_reset_reset_bridge_in_reset_reset                     : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                                   : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                               : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                      : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                                  : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                                     : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                               : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                            : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                        : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                               : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                           : out std_logic_vector(31 downto 0);                    -- readdata
			audio_avalon_audio_slave_address                          : out std_logic_vector(1 downto 0);                     -- address
			audio_avalon_audio_slave_write                            : out std_logic;                                        -- write
			audio_avalon_audio_slave_read                             : out std_logic;                                        -- read
			audio_avalon_audio_slave_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_avalon_audio_slave_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			audio_avalon_audio_slave_chipselect                       : out std_logic;                                        -- chipselect
			audio_and_video_config_avalon_av_config_slave_address     : out std_logic_vector(1 downto 0);                     -- address
			audio_and_video_config_avalon_av_config_slave_write       : out std_logic;                                        -- write
			audio_and_video_config_avalon_av_config_slave_read        : out std_logic;                                        -- read
			audio_and_video_config_avalon_av_config_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_and_video_config_avalon_av_config_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			audio_and_video_config_avalon_av_config_slave_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			audio_and_video_config_avalon_av_config_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_address                               : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                                 : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                                  : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable                            : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest                           : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess                           : out std_logic;                                        -- debugaccess
			DataFromAccMat_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			DataFromAccMat_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DataToAccMat_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			DataToAccMat_s1_write                                     : out std_logic;                                        -- write
			DataToAccMat_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DataToAccMat_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			DataToAccMat_s1_chipselect                                : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address                     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                       : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                        : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                  : out std_logic;                                        -- chipselect
			onchipmem_s1_address                                      : out std_logic_vector(15 downto 0);                    -- address
			onchipmem_s1_write                                        : out std_logic;                                        -- write
			onchipmem_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchipmem_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			onchipmem_s1_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			onchipmem_s1_chipselect                                   : out std_logic;                                        -- chipselect
			onchipmem_s1_clken                                        : out std_logic;                                        -- clken
			ps2_avalon_ps2_slave_address                              : out std_logic_vector(0 downto 0);                     -- address
			ps2_avalon_ps2_slave_write                                : out std_logic;                                        -- write
			ps2_avalon_ps2_slave_read                                 : out std_logic;                                        -- read
			ps2_avalon_ps2_slave_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ps2_avalon_ps2_slave_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			ps2_avalon_ps2_slave_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			ps2_avalon_ps2_slave_waitrequest                          : in  std_logic                     := 'X';             -- waitrequest
			ps2_avalon_ps2_slave_chipselect                           : out std_logic;                                        -- chipselect
			sysid_control_slave_address                               : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer0_s1_address                                         : out std_logic_vector(2 downto 0);                     -- address
			timer0_s1_write                                           : out std_logic;                                        -- write
			timer0_s1_readdata                                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer0_s1_writedata                                       : out std_logic_vector(15 downto 0);                    -- writedata
			timer0_s1_chipselect                                      : out std_logic;                                        -- chipselect
			timer1_s1_address                                         : out std_logic_vector(2 downto 0);                     -- address
			timer1_s1_write                                           : out std_logic;                                        -- write
			timer1_s1_readdata                                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer1_s1_writedata                                       : out std_logic_vector(15 downto 0);                    -- writedata
			timer1_s1_chipselect                                      : out std_logic;                                        -- chipselect
			ToggleAccMat_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			ToggleAccMat_s1_write                                     : out std_logic;                                        -- write
			ToggleAccMat_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ToggleAccMat_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			ToggleAccMat_s1_chipselect                                : out std_logic                                         -- chipselect
		);
	end component CodecAudio_mm_interconnect_0;

	component CodecAudio_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component CodecAudio_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component codecaudio_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component codecaudio_rst_controller;

	component codecaudio_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component codecaudio_rst_controller_001;

	signal dac_pll_audio_clk_clk                                                       : std_logic;                     -- dac_pll:audio_clk_clk -> [audio:clk, irq_synchronizer:receiver_clk, mm_interconnect_0:dac_pll_audio_clk_clk, rst_controller_001:clk]
	signal pll_0_outclk0_clk                                                           : std_logic;                     -- pll_0:outclk_0 -> [DataFromAccMat:clk, DataToAccMat:clk, ToggleAccMat:clk, audio_and_video_config:clk, cpu:clk, dac_pll:ref_clk_clk, dacchip_pll:ref_clk_clk, irq_mapper:clk, irq_synchronizer:sender_clk, jtag_uart_0:clk, mm_interconnect_0:pll_0_outclk0_clk, onchipmem:clk, ps2:clk, rst_controller:clk, sysid:clock, timer0:clk, timer1:clk]
	signal cpu_data_master_readdata                                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                                 : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                                 : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                                     : std_logic_vector(19 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                                  : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                                        : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                                       : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                                   : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                          : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                              : std_logic_vector(19 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                                 : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal mm_interconnect_0_audio_avalon_audio_slave_chipselect                       : std_logic;                     -- mm_interconnect_0:audio_avalon_audio_slave_chipselect -> audio:chipselect
	signal mm_interconnect_0_audio_avalon_audio_slave_readdata                         : std_logic_vector(31 downto 0); -- audio:readdata -> mm_interconnect_0:audio_avalon_audio_slave_readdata
	signal mm_interconnect_0_audio_avalon_audio_slave_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_avalon_audio_slave_address -> audio:address
	signal mm_interconnect_0_audio_avalon_audio_slave_read                             : std_logic;                     -- mm_interconnect_0:audio_avalon_audio_slave_read -> audio:read
	signal mm_interconnect_0_audio_avalon_audio_slave_write                            : std_logic;                     -- mm_interconnect_0:audio_avalon_audio_slave_write -> audio:write
	signal mm_interconnect_0_audio_avalon_audio_slave_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_avalon_audio_slave_writedata -> audio:writedata
	signal mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_readdata    : std_logic_vector(31 downto 0); -- audio_and_video_config:readdata -> mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_readdata
	signal mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_waitrequest : std_logic;                     -- audio_and_video_config:waitrequest -> mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_waitrequest
	signal mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_address     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_address -> audio_and_video_config:address
	signal mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_read        : std_logic;                     -- mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_read -> audio_and_video_config:read
	signal mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_byteenable -> audio_and_video_config:byteenable
	signal mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_write       : std_logic;                     -- mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_write -> audio_and_video_config:write
	signal mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_writedata -> audio_and_video_config:writedata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect                  : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata                    : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest                 : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                        : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write                       : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_ps2_avalon_ps2_slave_chipselect                           : std_logic;                     -- mm_interconnect_0:ps2_avalon_ps2_slave_chipselect -> ps2:chipselect
	signal mm_interconnect_0_ps2_avalon_ps2_slave_readdata                             : std_logic_vector(31 downto 0); -- ps2:readdata -> mm_interconnect_0:ps2_avalon_ps2_slave_readdata
	signal mm_interconnect_0_ps2_avalon_ps2_slave_waitrequest                          : std_logic;                     -- ps2:waitrequest -> mm_interconnect_0:ps2_avalon_ps2_slave_waitrequest
	signal mm_interconnect_0_ps2_avalon_ps2_slave_address                              : std_logic_vector(0 downto 0);  -- mm_interconnect_0:ps2_avalon_ps2_slave_address -> ps2:address
	signal mm_interconnect_0_ps2_avalon_ps2_slave_read                                 : std_logic;                     -- mm_interconnect_0:ps2_avalon_ps2_slave_read -> ps2:read
	signal mm_interconnect_0_ps2_avalon_ps2_slave_byteenable                           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ps2_avalon_ps2_slave_byteenable -> ps2:byteenable
	signal mm_interconnect_0_ps2_avalon_ps2_slave_write                                : std_logic;                     -- mm_interconnect_0:ps2_avalon_ps2_slave_write -> ps2:write
	signal mm_interconnect_0_ps2_avalon_ps2_slave_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:ps2_avalon_ps2_slave_writedata -> ps2:writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                              : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                               : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                              : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                           : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                           : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                               : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                                  : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                                 : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_onchipmem_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:onchipmem_s1_chipselect -> onchipmem:chipselect
	signal mm_interconnect_0_onchipmem_s1_readdata                                     : std_logic_vector(31 downto 0); -- onchipmem:readdata -> mm_interconnect_0:onchipmem_s1_readdata
	signal mm_interconnect_0_onchipmem_s1_address                                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:onchipmem_s1_address -> onchipmem:address
	signal mm_interconnect_0_onchipmem_s1_byteenable                                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchipmem_s1_byteenable -> onchipmem:byteenable
	signal mm_interconnect_0_onchipmem_s1_write                                        : std_logic;                     -- mm_interconnect_0:onchipmem_s1_write -> onchipmem:write
	signal mm_interconnect_0_onchipmem_s1_writedata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchipmem_s1_writedata -> onchipmem:writedata
	signal mm_interconnect_0_onchipmem_s1_clken                                        : std_logic;                     -- mm_interconnect_0:onchipmem_s1_clken -> onchipmem:clken
	signal mm_interconnect_0_timer0_s1_chipselect                                      : std_logic;                     -- mm_interconnect_0:timer0_s1_chipselect -> timer0:chipselect
	signal mm_interconnect_0_timer0_s1_readdata                                        : std_logic_vector(15 downto 0); -- timer0:readdata -> mm_interconnect_0:timer0_s1_readdata
	signal mm_interconnect_0_timer0_s1_address                                         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer0_s1_address -> timer0:address
	signal mm_interconnect_0_timer0_s1_write                                           : std_logic;                     -- mm_interconnect_0:timer0_s1_write -> mm_interconnect_0_timer0_s1_write:in
	signal mm_interconnect_0_timer0_s1_writedata                                       : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer0_s1_writedata -> timer0:writedata
	signal mm_interconnect_0_timer1_s1_chipselect                                      : std_logic;                     -- mm_interconnect_0:timer1_s1_chipselect -> timer1:chipselect
	signal mm_interconnect_0_timer1_s1_readdata                                        : std_logic_vector(15 downto 0); -- timer1:readdata -> mm_interconnect_0:timer1_s1_readdata
	signal mm_interconnect_0_timer1_s1_address                                         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer1_s1_address -> timer1:address
	signal mm_interconnect_0_timer1_s1_write                                           : std_logic;                     -- mm_interconnect_0:timer1_s1_write -> mm_interconnect_0_timer1_s1_write:in
	signal mm_interconnect_0_timer1_s1_writedata                                       : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer1_s1_writedata -> timer1:writedata
	signal mm_interconnect_0_toggleaccmat_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:ToggleAccMat_s1_chipselect -> ToggleAccMat:chipselect
	signal mm_interconnect_0_toggleaccmat_s1_readdata                                  : std_logic_vector(31 downto 0); -- ToggleAccMat:readdata -> mm_interconnect_0:ToggleAccMat_s1_readdata
	signal mm_interconnect_0_toggleaccmat_s1_address                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ToggleAccMat_s1_address -> ToggleAccMat:address
	signal mm_interconnect_0_toggleaccmat_s1_write                                     : std_logic;                     -- mm_interconnect_0:ToggleAccMat_s1_write -> mm_interconnect_0_toggleaccmat_s1_write:in
	signal mm_interconnect_0_toggleaccmat_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:ToggleAccMat_s1_writedata -> ToggleAccMat:writedata
	signal mm_interconnect_0_datatoaccmat_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:DataToAccMat_s1_chipselect -> DataToAccMat:chipselect
	signal mm_interconnect_0_datatoaccmat_s1_readdata                                  : std_logic_vector(31 downto 0); -- DataToAccMat:readdata -> mm_interconnect_0:DataToAccMat_s1_readdata
	signal mm_interconnect_0_datatoaccmat_s1_address                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:DataToAccMat_s1_address -> DataToAccMat:address
	signal mm_interconnect_0_datatoaccmat_s1_write                                     : std_logic;                     -- mm_interconnect_0:DataToAccMat_s1_write -> mm_interconnect_0_datatoaccmat_s1_write:in
	signal mm_interconnect_0_datatoaccmat_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:DataToAccMat_s1_writedata -> DataToAccMat:writedata
	signal mm_interconnect_0_datafromaccmat_s1_readdata                                : std_logic_vector(31 downto 0); -- DataFromAccMat:readdata -> mm_interconnect_0:DataFromAccMat_s1_readdata
	signal mm_interconnect_0_datafromaccmat_s1_address                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:DataFromAccMat_s1_address -> DataFromAccMat:address
	signal irq_mapper_receiver0_irq                                                    : std_logic;                     -- ps2:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver2_irq                                                    : std_logic;                     -- timer0:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                    : std_logic;                     -- timer1:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                                    : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver4_irq
	signal cpu_irq_irq                                                                 : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal irq_mapper_receiver1_irq                                                    : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	signal irq_synchronizer_receiver_irq                                               : std_logic_vector(0 downto 0);  -- audio:irq -> irq_synchronizer:receiver_irq
	signal rst_controller_reset_out_reset                                              : std_logic;                     -- rst_controller:reset_out -> [audio_and_video_config:reset, irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchipmem:reset, ps2:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                          : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, onchipmem:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                                          : std_logic;                     -- rst_controller_001:reset_out -> [audio:reset, irq_synchronizer:receiver_reset, mm_interconnect_0:audio_reset_reset_bridge_in_reset_reset]
	signal dac_pll_reset_source_reset                                                  : std_logic;                     -- dac_pll:reset_source_reset -> rst_controller_001:reset_in0
	signal reset_reset_n_ports_inv                                                     : std_logic;                     -- reset_reset_n:inv -> [dac_pll:ref_reset_reset, dacchip_pll:ref_reset_reset, pll_0:rst, rst_controller:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv              : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv             : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_timer0_s1_write_ports_inv                                 : std_logic;                     -- mm_interconnect_0_timer0_s1_write:inv -> timer0:write_n
	signal mm_interconnect_0_timer1_s1_write_ports_inv                                 : std_logic;                     -- mm_interconnect_0_timer1_s1_write:inv -> timer1:write_n
	signal mm_interconnect_0_toggleaccmat_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_toggleaccmat_s1_write:inv -> ToggleAccMat:write_n
	signal mm_interconnect_0_datatoaccmat_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_datatoaccmat_s1_write:inv -> DataToAccMat:write_n
	signal rst_controller_reset_out_reset_ports_inv                                    : std_logic;                     -- rst_controller_reset_out_reset:inv -> [DataFromAccMat:reset_n, DataToAccMat:reset_n, ToggleAccMat:reset_n, cpu:reset_n, jtag_uart_0:rst_n, sysid:reset_n, timer0:reset_n, timer1:reset_n]

begin

	datafromaccmat : component CodecAudio_DataFromAccMat
		port map (
			clk      => pll_0_outclk0_clk,                            --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address  => mm_interconnect_0_datafromaccmat_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_datafromaccmat_s1_readdata, --                    .readdata
			in_port  => datafromaccmat_i_export                       -- external_connection.export
		);

	datatoaccmat : component CodecAudio_DataToAccMat
		port map (
			clk        => pll_0_outclk0_clk,                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_datatoaccmat_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_datatoaccmat_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_datatoaccmat_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_datatoaccmat_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_datatoaccmat_s1_readdata,        --                    .readdata
			out_port   => datatoaccmat_o_export                              -- external_connection.export
		);

	toggleaccmat : component CodecAudio_ToggleAccMat
		port map (
			clk        => pll_0_outclk0_clk,                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_toggleaccmat_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_toggleaccmat_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_toggleaccmat_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_toggleaccmat_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_toggleaccmat_s1_readdata,        --                    .readdata
			in_port    => toggleaccmat_i_export                              -- external_connection.export
		);

	audio : component CodecAudio_audio
		port map (
			clk         => dac_pll_audio_clk_clk,                                 --                clk.clk
			reset       => rst_controller_001_reset_out_reset,                    --              reset.reset
			address     => mm_interconnect_0_audio_avalon_audio_slave_address,    -- avalon_audio_slave.address
			chipselect  => mm_interconnect_0_audio_avalon_audio_slave_chipselect, --                   .chipselect
			read        => mm_interconnect_0_audio_avalon_audio_slave_read,       --                   .read
			write       => mm_interconnect_0_audio_avalon_audio_slave_write,      --                   .write
			writedata   => mm_interconnect_0_audio_avalon_audio_slave_writedata,  --                   .writedata
			readdata    => mm_interconnect_0_audio_avalon_audio_slave_readdata,   --                   .readdata
			irq         => irq_synchronizer_receiver_irq(0),                      --          interrupt.irq
			AUD_BCLK    => audio_o_BCLK,                                          -- external_interface.export
			AUD_DACDAT  => audio_o_DACDAT,                                        --                   .export
			AUD_DACLRCK => audio_o_DACLRCK                                        --                   .export
		);

	audio_and_video_config : component CodecAudio_audio_and_video_config
		port map (
			clk         => pll_0_outclk0_clk,                                                           --                    clk.clk
			reset       => rst_controller_reset_out_reset,                                              --                  reset.reset
			address     => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_address,     -- avalon_av_config_slave.address
			byteenable  => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_byteenable,  --                       .byteenable
			read        => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_read,        --                       .read
			write       => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_write,       --                       .write
			writedata   => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_writedata,   --                       .writedata
			readdata    => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_readdata,    --                       .readdata
			waitrequest => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_waitrequest, --                       .waitrequest
			I2C_SDAT    => audio_i2c_o_SDAT,                                                            --     external_interface.export
			I2C_SCLK    => audio_i2c_o_SCLK                                                             --                       .export
		);

	cpu : component CodecAudio_cpu
		port map (
			clk                                 => pll_0_outclk0_clk,                                 --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                              --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	dac_pll : component CodecAudio_dac_pll
		port map (
			ref_clk_clk        => pll_0_outclk0_clk,          --      ref_clk.clk
			ref_reset_reset    => reset_reset_n_ports_inv,    --    ref_reset.reset
			audio_clk_clk      => dac_pll_audio_clk_clk,      --    audio_clk.clk
			reset_source_reset => dac_pll_reset_source_reset  -- reset_source.reset
		);

	dacchip_pll : component CodecAudio_dac_pll
		port map (
			ref_clk_clk        => pll_0_outclk0_clk,         --      ref_clk.clk
			ref_reset_reset    => reset_reset_n_ports_inv,   --    ref_reset.reset
			audio_clk_clk      => dacchip_pll_audio_clk_clk, --    audio_clk.clk
			reset_source_reset => open                       -- reset_source.reset
		);

	jtag_uart_0 : component CodecAudio_jtag_uart_0
		port map (
			clk            => pll_0_outclk0_clk,                                               --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver4_irq                                         --               irq.irq
		);

	onchipmem : component CodecAudio_onchipmem
		port map (
			clk        => pll_0_outclk0_clk,                         --   clk1.clk
			address    => mm_interconnect_0_onchipmem_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchipmem_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchipmem_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchipmem_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchipmem_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchipmem_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchipmem_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,            -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req         --       .reset_req
		);

	pll_0 : component CodecAudio_pll_0
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_0_outclk0_clk,       -- outclk0.clk
			locked   => pll_0_locked_export      --  locked.export
		);

	ps2 : component CodecAudio_ps2
		port map (
			clk         => pll_0_outclk0_clk,                                  --                clk.clk
			reset       => rst_controller_reset_out_reset,                     --              reset.reset
			address     => mm_interconnect_0_ps2_avalon_ps2_slave_address(0),  --   avalon_ps2_slave.address
			chipselect  => mm_interconnect_0_ps2_avalon_ps2_slave_chipselect,  --                   .chipselect
			byteenable  => mm_interconnect_0_ps2_avalon_ps2_slave_byteenable,  --                   .byteenable
			read        => mm_interconnect_0_ps2_avalon_ps2_slave_read,        --                   .read
			write       => mm_interconnect_0_ps2_avalon_ps2_slave_write,       --                   .write
			writedata   => mm_interconnect_0_ps2_avalon_ps2_slave_writedata,   --                   .writedata
			readdata    => mm_interconnect_0_ps2_avalon_ps2_slave_readdata,    --                   .readdata
			waitrequest => mm_interconnect_0_ps2_avalon_ps2_slave_waitrequest, --                   .waitrequest
			irq         => irq_mapper_receiver0_irq,                           --          interrupt.irq
			PS2_CLK     => ps2_o_CLK,                                          -- external_interface.export
			PS2_DAT     => ps2_o_DAT                                           --                   .export
		);

	sysid : component CodecAudio_sysid
		port map (
			clock    => pll_0_outclk0_clk,                                --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	timer0 : component CodecAudio_timer0
		port map (
			clk        => pll_0_outclk0_clk,                           --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    -- reset.reset_n
			address    => mm_interconnect_0_timer0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                     --   irq.irq
		);

	timer1 : component CodecAudio_timer1
		port map (
			clk        => pll_0_outclk0_clk,                           --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    -- reset.reset_n
			address    => mm_interconnect_0_timer1_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer1_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer1_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer1_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer1_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver3_irq                     --   irq.irq
		);

	mm_interconnect_0 : component CodecAudio_mm_interconnect_0
		port map (
			dac_pll_audio_clk_clk                                     => dac_pll_audio_clk_clk,                                                       --                             dac_pll_audio_clk.clk
			pll_0_outclk0_clk                                         => pll_0_outclk0_clk,                                                           --                                 pll_0_outclk0.clk
			audio_reset_reset_bridge_in_reset_reset                   => rst_controller_001_reset_out_reset,                                          --             audio_reset_reset_bridge_in_reset.reset
			cpu_reset_reset_bridge_in_reset_reset                     => rst_controller_reset_out_reset,                                              --               cpu_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                                   => cpu_data_master_address,                                                     --                               cpu_data_master.address
			cpu_data_master_waitrequest                               => cpu_data_master_waitrequest,                                                 --                                              .waitrequest
			cpu_data_master_byteenable                                => cpu_data_master_byteenable,                                                  --                                              .byteenable
			cpu_data_master_read                                      => cpu_data_master_read,                                                        --                                              .read
			cpu_data_master_readdata                                  => cpu_data_master_readdata,                                                    --                                              .readdata
			cpu_data_master_write                                     => cpu_data_master_write,                                                       --                                              .write
			cpu_data_master_writedata                                 => cpu_data_master_writedata,                                                   --                                              .writedata
			cpu_data_master_debugaccess                               => cpu_data_master_debugaccess,                                                 --                                              .debugaccess
			cpu_instruction_master_address                            => cpu_instruction_master_address,                                              --                        cpu_instruction_master.address
			cpu_instruction_master_waitrequest                        => cpu_instruction_master_waitrequest,                                          --                                              .waitrequest
			cpu_instruction_master_read                               => cpu_instruction_master_read,                                                 --                                              .read
			cpu_instruction_master_readdata                           => cpu_instruction_master_readdata,                                             --                                              .readdata
			audio_avalon_audio_slave_address                          => mm_interconnect_0_audio_avalon_audio_slave_address,                          --                      audio_avalon_audio_slave.address
			audio_avalon_audio_slave_write                            => mm_interconnect_0_audio_avalon_audio_slave_write,                            --                                              .write
			audio_avalon_audio_slave_read                             => mm_interconnect_0_audio_avalon_audio_slave_read,                             --                                              .read
			audio_avalon_audio_slave_readdata                         => mm_interconnect_0_audio_avalon_audio_slave_readdata,                         --                                              .readdata
			audio_avalon_audio_slave_writedata                        => mm_interconnect_0_audio_avalon_audio_slave_writedata,                        --                                              .writedata
			audio_avalon_audio_slave_chipselect                       => mm_interconnect_0_audio_avalon_audio_slave_chipselect,                       --                                              .chipselect
			audio_and_video_config_avalon_av_config_slave_address     => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_address,     -- audio_and_video_config_avalon_av_config_slave.address
			audio_and_video_config_avalon_av_config_slave_write       => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_write,       --                                              .write
			audio_and_video_config_avalon_av_config_slave_read        => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_read,        --                                              .read
			audio_and_video_config_avalon_av_config_slave_readdata    => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_readdata,    --                                              .readdata
			audio_and_video_config_avalon_av_config_slave_writedata   => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_writedata,   --                                              .writedata
			audio_and_video_config_avalon_av_config_slave_byteenable  => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_byteenable,  --                                              .byteenable
			audio_and_video_config_avalon_av_config_slave_waitrequest => mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_waitrequest, --                                              .waitrequest
			cpu_debug_mem_slave_address                               => mm_interconnect_0_cpu_debug_mem_slave_address,                               --                           cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                                 => mm_interconnect_0_cpu_debug_mem_slave_write,                                 --                                              .write
			cpu_debug_mem_slave_read                                  => mm_interconnect_0_cpu_debug_mem_slave_read,                                  --                                              .read
			cpu_debug_mem_slave_readdata                              => mm_interconnect_0_cpu_debug_mem_slave_readdata,                              --                                              .readdata
			cpu_debug_mem_slave_writedata                             => mm_interconnect_0_cpu_debug_mem_slave_writedata,                             --                                              .writedata
			cpu_debug_mem_slave_byteenable                            => mm_interconnect_0_cpu_debug_mem_slave_byteenable,                            --                                              .byteenable
			cpu_debug_mem_slave_waitrequest                           => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,                           --                                              .waitrequest
			cpu_debug_mem_slave_debugaccess                           => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,                           --                                              .debugaccess
			DataFromAccMat_s1_address                                 => mm_interconnect_0_datafromaccmat_s1_address,                                 --                             DataFromAccMat_s1.address
			DataFromAccMat_s1_readdata                                => mm_interconnect_0_datafromaccmat_s1_readdata,                                --                                              .readdata
			DataToAccMat_s1_address                                   => mm_interconnect_0_datatoaccmat_s1_address,                                   --                               DataToAccMat_s1.address
			DataToAccMat_s1_write                                     => mm_interconnect_0_datatoaccmat_s1_write,                                     --                                              .write
			DataToAccMat_s1_readdata                                  => mm_interconnect_0_datatoaccmat_s1_readdata,                                  --                                              .readdata
			DataToAccMat_s1_writedata                                 => mm_interconnect_0_datatoaccmat_s1_writedata,                                 --                                              .writedata
			DataToAccMat_s1_chipselect                                => mm_interconnect_0_datatoaccmat_s1_chipselect,                                --                                              .chipselect
			jtag_uart_0_avalon_jtag_slave_address                     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,                     --                 jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,                       --                                              .write
			jtag_uart_0_avalon_jtag_slave_read                        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,                        --                                              .read
			jtag_uart_0_avalon_jtag_slave_readdata                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,                    --                                              .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,                   --                                              .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                 => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,                 --                                              .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,                  --                                              .chipselect
			onchipmem_s1_address                                      => mm_interconnect_0_onchipmem_s1_address,                                      --                                  onchipmem_s1.address
			onchipmem_s1_write                                        => mm_interconnect_0_onchipmem_s1_write,                                        --                                              .write
			onchipmem_s1_readdata                                     => mm_interconnect_0_onchipmem_s1_readdata,                                     --                                              .readdata
			onchipmem_s1_writedata                                    => mm_interconnect_0_onchipmem_s1_writedata,                                    --                                              .writedata
			onchipmem_s1_byteenable                                   => mm_interconnect_0_onchipmem_s1_byteenable,                                   --                                              .byteenable
			onchipmem_s1_chipselect                                   => mm_interconnect_0_onchipmem_s1_chipselect,                                   --                                              .chipselect
			onchipmem_s1_clken                                        => mm_interconnect_0_onchipmem_s1_clken,                                        --                                              .clken
			ps2_avalon_ps2_slave_address                              => mm_interconnect_0_ps2_avalon_ps2_slave_address,                              --                          ps2_avalon_ps2_slave.address
			ps2_avalon_ps2_slave_write                                => mm_interconnect_0_ps2_avalon_ps2_slave_write,                                --                                              .write
			ps2_avalon_ps2_slave_read                                 => mm_interconnect_0_ps2_avalon_ps2_slave_read,                                 --                                              .read
			ps2_avalon_ps2_slave_readdata                             => mm_interconnect_0_ps2_avalon_ps2_slave_readdata,                             --                                              .readdata
			ps2_avalon_ps2_slave_writedata                            => mm_interconnect_0_ps2_avalon_ps2_slave_writedata,                            --                                              .writedata
			ps2_avalon_ps2_slave_byteenable                           => mm_interconnect_0_ps2_avalon_ps2_slave_byteenable,                           --                                              .byteenable
			ps2_avalon_ps2_slave_waitrequest                          => mm_interconnect_0_ps2_avalon_ps2_slave_waitrequest,                          --                                              .waitrequest
			ps2_avalon_ps2_slave_chipselect                           => mm_interconnect_0_ps2_avalon_ps2_slave_chipselect,                           --                                              .chipselect
			sysid_control_slave_address                               => mm_interconnect_0_sysid_control_slave_address,                               --                           sysid_control_slave.address
			sysid_control_slave_readdata                              => mm_interconnect_0_sysid_control_slave_readdata,                              --                                              .readdata
			timer0_s1_address                                         => mm_interconnect_0_timer0_s1_address,                                         --                                     timer0_s1.address
			timer0_s1_write                                           => mm_interconnect_0_timer0_s1_write,                                           --                                              .write
			timer0_s1_readdata                                        => mm_interconnect_0_timer0_s1_readdata,                                        --                                              .readdata
			timer0_s1_writedata                                       => mm_interconnect_0_timer0_s1_writedata,                                       --                                              .writedata
			timer0_s1_chipselect                                      => mm_interconnect_0_timer0_s1_chipselect,                                      --                                              .chipselect
			timer1_s1_address                                         => mm_interconnect_0_timer1_s1_address,                                         --                                     timer1_s1.address
			timer1_s1_write                                           => mm_interconnect_0_timer1_s1_write,                                           --                                              .write
			timer1_s1_readdata                                        => mm_interconnect_0_timer1_s1_readdata,                                        --                                              .readdata
			timer1_s1_writedata                                       => mm_interconnect_0_timer1_s1_writedata,                                       --                                              .writedata
			timer1_s1_chipselect                                      => mm_interconnect_0_timer1_s1_chipselect,                                      --                                              .chipselect
			ToggleAccMat_s1_address                                   => mm_interconnect_0_toggleaccmat_s1_address,                                   --                               ToggleAccMat_s1.address
			ToggleAccMat_s1_write                                     => mm_interconnect_0_toggleaccmat_s1_write,                                     --                                              .write
			ToggleAccMat_s1_readdata                                  => mm_interconnect_0_toggleaccmat_s1_readdata,                                  --                                              .readdata
			ToggleAccMat_s1_writedata                                 => mm_interconnect_0_toggleaccmat_s1_writedata,                                 --                                              .writedata
			ToggleAccMat_s1_chipselect                                => mm_interconnect_0_toggleaccmat_s1_chipselect                                 --                                              .chipselect
		);

	irq_mapper : component CodecAudio_irq_mapper
		port map (
			clk           => pll_0_outclk0_clk,              --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,       -- receiver4.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => dac_pll_audio_clk_clk,              --       receiver_clk.clk
			sender_clk     => pll_0_outclk0_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_001_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_reset_out_reset,     --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver1_irq            --             sender.irq
		);

	rst_controller : component codecaudio_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => pll_0_outclk0_clk,                  --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component codecaudio_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => dac_pll_reset_source_reset,         -- reset_in0.reset
			clk            => dac_pll_audio_clk_clk,              --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_timer0_s1_write_ports_inv <= not mm_interconnect_0_timer0_s1_write;

	mm_interconnect_0_timer1_s1_write_ports_inv <= not mm_interconnect_0_timer1_s1_write;

	mm_interconnect_0_toggleaccmat_s1_write_ports_inv <= not mm_interconnect_0_toggleaccmat_s1_write;

	mm_interconnect_0_datatoaccmat_s1_write_ports_inv <= not mm_interconnect_0_datatoaccmat_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of CodecAudio
