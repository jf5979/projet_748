// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ywDRFLKJKUG8cnHcgGtV0evrGJro3RXg6RPWf1LW8Ug2gvukxC2Bzfw+2gbwtau39tkqe4DMptda
73h0TnFYHjuxrR3CL1B8zTzH/V0X/5rT8nmze9mIz7Xlcq/bBNHIK4sfRZt2GKZv3ggDy/3RvwI4
lhWXD58hUAP9aorEUVwMwVGMnD3tZlPZu1Ug+2hoNhp3l9qUCXBKqoBAwIi15aPyZD7TqHUc1HDE
gruImTJZ6kEeNjBFENeDGCqkk5TjneggzbfanoyNSECyh76q4kd3hIM3dOHHnIL2QlTXPWP74Yrn
Ynyv8gEZfyKOdeqiFZ80JbejCB6S5aLq2BAbzw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17376)
Nf5yoh24xxjx7j78ukSo2/D5mF9sG5LdgrhiBSBr5TjYcvPtDmwrBGLXyx7oxXV7atZn5Xh6fg1p
yZ6Yb9Zqb4vU9LLUtML/mDTwBrkuv8wct+aPesjphlNobcekS2k6vuSVZLMEzxJ2erabWWU36bsN
acixvJyzBUmNiLQGb1eugpEOU8AMvRfThbfRAh3/YU4juFsoB9OMHNqMoZ1oguveRp9wejM57BSi
7qksf8/6eUQgTmz/Vw+ts8Ow0mL4yelhUePXjkLkjJqq+9pM+eXl0DPmAjFEFekl+35MqLfumR3m
BBNb18AdQc1VcVaKEsDCVzA7nORAxG8nNxh+53n6hcebJuXSfCVnY/1qKy9yBPOvv08G97j/jN3+
7NOcNWYw9Ei/Brk/5tzFtDVBnZ86GDRLRQl62PFpJ40DyOjKM5tEVRFc+6+GgyQQ3AfdGk5DWXri
LHv3zkPm8kkWjXxovLL75w2U7aO1IOFt4iiIBewH3FgG/ocQ6hAmtkV4PcveD5pd+6d2f3d2C8Jx
1GF3R1hL6qbtyE6NN+EQE/ecCNHevcEp0lmIlxuV/rUdgvRw9gKlIM3L1BnP9czc4pA+vNX9/MEW
kGsH0vQDA1WrSJOEnUX0wKsPoDzyaL8rfPzaUwUdFHeb8ENi7V7/PAqar0MhfQ+14wgSBCvQHruQ
5eHPO+J7TZp4dSukGnK418oL2nOIVBCOXvJ5lBZzsDxnvfM3Dvh6PdLe7XCFTWsSaRMCQDWp4Ctd
I8IxfzqQx0NAQWNIqkhPCOr8ZSgkFxI4j7QBB3DMy0qecOhPrp9YVkEbDY0s9mDMbeZ1hfKlibot
C5q8ZsjH6EZ1LZzjnsIfdQtYJ3oq97gSamRrc+woeO2mqvH0DyS/xkNShRI2tQxpZzV9K5AeBAkr
rEiyDuZw3hAJ4dz9/SgVN9AqoXMzV5PSJXpWihoixO0CAYz+o8GOD5WEgVY7EJwJGM5Yrwsf8WCp
AcS435GbU0OUgpMeMcs9SGR88Cr5pYmPoo+ulUVQk1wORokCU+NPtDJrdUVlYDiJhT43CWP0Iu6x
HUXc//Q/8rxBcT0StUvVcrF1fBmQFAwa+faDww0acSfljJ7C3ufX6/YPCdS9ef3jGu/zT5TtR109
O3jXBmsxgUZA0RayadCHNIGwVqKC9qO0Bx8SV1B6yQ3H8KMBIEsoun3fggnk0LyZb1l28ASAJTHe
oZzIIfcRavbGs6Yv6mtoVmAabYyeitOqOq2I5P5iqHllZS0qKj2YjEnItrPTMjjlL12jhIdvgjqf
VNIqWkaGYVSYLrGjPHt+l7drTVUTm3QEgV2mX+voBmGJrFVhcaU9618LRFWDuNWpJ9HdptINKPii
C80DFv+muOuG1FAQmNgUcfp2qsLNJi7DKWLL+Nj6nmszdhT5UPVOYmP2IMeh6UayPcORUNZDJIOh
wMQdYtVsCenHRB53wYBMQk0nxkazeu+x7Bwv9dbm5RFvCGcbC3s9aJtniZrhiA4Sq73EAla6CcAR
/hf6oJ7MmjRacdz9Cl0jIzHi9wSdnrXfwuU8RbEBi6rKAXfA1Mk25bgpFNuR5gYkpf2YapiAt3g4
Zrmbdr8sn1KkZxKj2Ie0hi4beP+CQC3Dd8JZu0BFj2ZYlGF0AMgteK1sLoF183Vz0QzCgAEeZYEs
ioiTm7PsC69YkdGiqkH4uddWNOWNo/Gs6aKLkyS+zq7LqvLASktryc35K3KVQO5SyF4NCdBAbEpR
y646v/s9oi8LmdeDAFsLaCttIcPsVAl2Kn0FYuSv9PRt4iSyMmNL+iCriQat3XDsOaw8WQmhKQ6p
d3p3OM7xaaUNFF0kG3XpD4iBqpCtuuo5T/YpW5iDT4AXVyTHNOrvDwZe8Z3mZTr/crpwHUklFbsk
63Xc45Qe3ydV5hxqpIJsmCHp3xGjwrsPiBPmhabKPIk8Cmje/2joOpRV6N+6fObKjRlHL06sOczj
t4GRDXI9fJe/IsxehSxlyaIe3PzLU2TjVVmvWqsIB+bonA7oPOaoejxkOsCGWpz63zIgB69Kooym
rIrasKBZ7mkw0319cLyqQVak6btd8JV5QRN/EUjfU8u2qdB1mp7y6+3jBZxuzCpfMfbjQ3NQ8ALy
BiIlTmn+X7Fx9uZXGLPBHq+qazbuHcIlb7QC5FY8uuG09bROe0FqszdP2iW86czU2WyUeCTxrkpD
Hf8FPrpQyiIEydyj3PX2T1cn+kXYdjGbziHmS9MOTYYhlK5DcddJeVjb0aeaLGdGF0xiZGDS7HxI
c3XtnNw7DBHeXnM7Te63LWOx1MbIjaNoLkZHj3ST1oPfwnoYiVURwJKfVnH7F4Flf71TQIkO2wWu
DkNJmygqChsDMCKqHixiPDaivJkF1/r/UYM4W9WjeUkl5NC51LRZrBfyNkjaRRlD7bxl+uJoankG
WY98UgQdWvQpd2bQfTcNbRxBzaHY8Kci5zUcswxJ2bcKBTk7CY0/Vi+7TzkKpGTv0C1sHQi9H+He
J9W3V0ioOgF87d3eKe1+aSAKpkOoDlSLW/zuzjCF+2yaPwYJKSyoU1L13wSnzYPuFid0xk/IfZQM
lfgiHPzpYiw/fx4AW1WDMkJNKTPGTqPHM9PO08tujPiHjUnbpoSrZ1xxioj3Uu4Q1hjw3uHYstyz
CFhBCJ9V1BXUrs4csRVLnww3Twzn1r2Aaft5MHcvh2o2cr5k7QnBsCEDL5CgfkffguLu3u1UJgyq
/7lTdS3xypT+Z1AzHj/7jwVUsKbu78afz1qtvrz6hes1ygd2bKpfqhwn2ytCLTdXrBWB6sE6mVJV
By2riLDoQn/1JBYLA9yOqfp23fGhj2kWSeQUspudwBpzcTORwl8m/SbFaV8r6U1OCLPFFIWgY/33
VYnO2ArR6ypWCwOpOoyq4ZJb23dNPtlUhCGyoglLX8VHlq9jBFgCpRz7vsrpLnH+B7DY3hKoZiOn
BpCJim3hD0GwuPqQlHa6Nj73UR0t6jex4eOrCw+K59l0Gd/eDafOzCIHhtFj/Ni0j0TQUsZYn99L
Egnfcqg58yPIfNP7uiR55zZ5uxAFHgsTO+v4b8gkYlxp46wv3s22bOXVSa1FdAJALxC//5GrOkKN
qLQ0+Qxbsry9rqnmv8h03wAamraZg3OmsSSHlC/UN87Td3yq1OPnUaoiFy6bESqscTcrSCb1oUoL
BtbPo1pbaSicxnJUn8znChsPRd8zRZ9K0Wj1sZxLuO8y5hFGBxptGkBHKN8TFui7bXkqFjz5DY/6
NvLrKs0XJzVM7tED7zU6kMIY5CHKwsG3jzvO+SBAYAZg5Puo0DMMuXmeTpPk6aYWi7QlzzbvEJmo
u8NHCMM3WqxxEpxzI1y3cThC6IoRdLI+fxEJr44G1UxWn+y4xU8drrTSWJ9sRuuksQPoWvCT9zVo
vHodY6eTlSwIn/HYXRCY+JrFOikuq0DYUm9uHP/SYlTlbVd81N9OxuZjEYYq+wFFsZTShPY/JewA
V8t0c71X4nlqCV5MEY4m7CQVS8lyWIhJqXrsQa0Ss4uqyWzX2+wSp+5nJLy83nrlj4g30Q5MOCsy
eKjrr43p9zzE9FfPE9CbLxod0YkzkPgGgPYmNlKm6H10+oc5wKET6VmG4sDmYdBuX7BKVVYTrGX6
SMIz3Nrq/sn2O7HQB54Z3rIEC8inR9y2nMFG1E0GOAm8Osc+NHONL77Ip49e2W5tVHrdR3zaxKXf
AdJsIEQMUSqfX4VVCEJZ7ui79V9fTXwLYlXzwVMXohEVdiWjDmudX0FxcwDWIVBoF9BP+iWCRqrb
BgFjn1R7q5v1W0ctlKvt78cZrnS25l4CRlTjzf6vmlQrmQ6AjyvzSyizelOx/kCRwPpq8eixjbt3
eqjTm9MkOvbbO/74eeR5tU6WEYc7mByKHY72HKP2Wfr4Ro+BrwRyIVthNYdoz7p1CGvvpYJ1Ozd1
uUCN0QyDDq2X/RxRb4ZNSYhH27tMscxg1VO63HjI1bKMrrB3/x+GEiEupnxVIJGIGjFd+u4BPJAy
5Qv9lZs/QAfzCU/D4xjdLqxJKDD4cWZOD+swFyyYY/zJirzRbJFlBNl1xKpj0oZE39f4kgJ+HCe0
x9SKiPG3Aqudg/7+qk8O0yhKSzR64j5jwpQHrEs99jl2xlRBSlSS/+BMWOIJx3rmw/6Bv9leao3o
4jPyRzd1ihjBg6vxk3OZ8L0Jc8HL5aPo5wt+0Mlr8bGPATWmnUEYLpMWFxYCVf0d91Kyv0X8ND5H
h8fLQOsS3CF2h2ZTRGrZaXeBXmiOU5nklMgFZm2f6Ai7vc09iZh8MuranBagVTEOMrDIuUmVRJTz
AIooqg27rboz0Lnaox+9ggakpT0Zl7NKYAOW5/11B8X9sslxdu0tD2aU5CtHANmUHvztQCNA++Ub
mYcg1LjSh/tXcPz0aV4W5yGKK546/aZW/jdzPvI8YdiF4jRAzZAAAyGb/gwzRUhFrjyCUOwB013Z
HRdFcDBK9eZlNuokpT+0AZE768Qysr18b+GRXJB9DGi8AYRW+49RN1zyRYXZKOTWyGYHdQuNR8Fz
7rcDmjur3kiKruUvyWQdLsJfqujQiZOrf2lQQsjwUuvNrOFLGN6w5f0QgEG17tQQwjeDZePmboD4
ADneg6pvjh76KUb31mvyGSUNeg3U7hozclTIF+qmkEqB3t8h6Ojh0LXrfkwzyAypBjUzcWPzgHyN
iI1s3HvfUnE9UwQYf/1zosAFhQIGJW5jCXSMxl9BeV71gN0jOnhiCWeVXE++O5wEA/4v5lkCJBkC
qHLIjq899ArWK4nnD0pUDrq9Mhi5pmB3OrGBxUGy1zNs0IbfiQb/ClQ3pLjpjpJ+wJuI6e7rC7AP
VIfJdJ6OxhWXUYS20UcuXVN3rv0+8T0hxPC0FeDj4vmvmnIAYHKhm+waGxz9xVtn47aDbKggd0GE
cp2UTjqgt8ki11hdOL5r8KhK7cB5lcUmLXWsvdzrP5eHTYLQr6q/KxE3O4jFBp9Oxq//ve/g5AOZ
VdVI9kvJ9X8Bn6vJD+KKLxDUu6oTdpPheZxRFrAgBCprwJCN3BFQndNEFVXjvtG1PzdRiB/YMDkg
lOovN7hyhUtdAN6MS8jVa/E/BEG2kyES6cT/f4Z/DWYtNwlKyujvpyOOnm7zRqUQne0qDkfrhjeq
GRo0jQzuqr9a9vlZM4Ga/zQPw49BTrnb8c7jUjlDGb8ggaahWCmZjaUa6g8oiI8m88tgNj9KVenR
xZD+1nV3KAL7GV8kyCo5UrM30g39vn17rpwsdPkvSyTfJAj9xm7HjpH129EEo/9a8HKELz/QU++y
Q9FxxD0AeGSpBfIaPAxTCyv+0UVgBZqfMyxOVaq0AIDtLlKwayEFzkClr0xrGYjHUycL2GBlQVSk
GnrS4l+GmAhanNIIEg7SzcWUYhXhsETXXrXsZTg06lWmNPpDI8iBLjK1gZYyMUpq9F0PzEDy/sWE
4UMU4iiL3tSy2vQi0UEF0OPKCm9/wwOikrBmP2Pso9BB96cUjtNrOmht/nDzQVP53vY3CfNG51/S
+PhZv1YgLgZc0W2qSShQkisJvkg2EPSC+RhgOcdt14f6My8DRKKIcx7kxUDED+5LQR4y0MBhIAaD
sYcjncUx8gdCa3ik11TZHLo9aYlHLLATN8YLekTtnndfsJt3IaK7TqBjot2ep2prLaNBQY99Ooln
eXSEBth2fFI+uG/dZNwoGizLCzBUnWAyg7lxG2bFMYFvMkDxtc3SSQaSVSiSj7cZOyBbks7LE+d2
FUE564D2+WqA8dHhRVD99PPNloepoca/7H6YpAoLp+PBSQiGJI0vnMtJRVzs3oLeHSc+33pG4vyq
QQuAeGd/J6XbqZcgiP0ZXa58iqd9FFppALzScMNbwxfAGBTzMzDSWlNjaX6J2F5ug/yKz1IbcjPv
RzFhoJIxqAvOkKfgoOBmvyR4QeyQ74zRdVQ8LRN0eFpzl0ou5a6uxnt0H4mKFuisN7XqPjGPZLBc
A5YmBnirNY/yLZPNsDBbxn0nOxENn+2mX2wMUZeLbLhXM9fn5E+Nq7k15pRYpD/zXuubcIKH9wnW
1Hsr3Qsi/Las4bMNZNVEr0nmjdWRyJky1q9LpQkxXzrzghpUm1BiLUol+TirrEbS+qS7O2wHIb68
IhdfmOn/Q68fPvsOijDo6U4b3nZSD1MgfKNh3Enq8x71wiygInbQuSz15ZFyN7FloelEFRTbs+7J
AkWkHJnzK2ObYw6pYbVEEcsVv0h/GZZrjMRR20p+cy/9BLCACGPsehnohKx45ANtg8+sm5kvFJpY
fvqRf6NEUhsX34qLIuLTTFXkVOo7iN3o4wl/QM37u903QY0Is5iLdKYXunbGaSAbO6Q1U97fmziK
hBo/rTMWoRdZrVdp/zEURKsi8HBwEmdq52FKkIo4sdI4k1jE0Yi7bVSnPugcC/ZNDuE6NgZc+xa2
TweJMOb/6BOWeqGpKu0mYZ7M7zG8LNRzRqrUfw2y48aLlDOXtfGxSTXDHbpiTTGdrrVr72vyMymf
74iF0+eUpB15oH2BerUwzcytR6hlS8jhfmxwYW4lxhv8yhbd3wd+1+wY7jNMti7SxQmoy9lhRdp1
LKkcN9t/UkaaYchNbRHc7qH3pUGLbsVqvOAulO4t628hBmvZ63FTKB5yol2FXdXzedcSWpm67YH0
B+B5Hm58E0hzg5G7Z1t1bJNacKeqLpWHxwes0fJHYi1oQyqGXkBYF+1hwMk0/KbaFIGFcLrXE373
QM1BZbeGi4vyPZGp9uv1fXaPF2p8xiubo87Z4sQS7DCjgLQlk5UC0lQ7aGRksCF2Y8S5tpDcwM12
Jd1SIJ13Lf5GSpGmU7QMqcf4xVeslk8GjVZWYj09PwYpfuxFRfEHFU/+FkD7NkYsq2WboVaFMrrB
TTyd3kKNIJ/vqh1WqlMAxYB7p9FBC+ou1U4dT1cnPB7UvOBRDEI9bXB733ZYVv9dhV9KKwKVWnWA
WN/xp8Q0SA3cONeYX9Vye+ylUdGYljtyM5WuQ8hsUwlYBgdXhuvJUqdqch/pWOxRSQDftdlFwBqJ
kBN07YIuoZIW2/305x/+CiZXnMM3bfF3CmmJYecsz7tbQuyOX+MUXI61cLmphYCmQOHdeeazIedo
+kCfQR44d3JReNJxFMN47AHol9C4Fo6D9KJE9lIqJBFFFYbHF2GJUiWe/9Y01p3swS1fjYb1+RN5
MK9rHFe9XOsU0ESshwIBk0SO4W/DlRzNWIIrtR4oJenKPl9OceSDJ7a5rRs88wZGg6fRDrcQv5Ct
il1we86Gt1WEy0rJQIlwFGlsEY1FqVpssxi/kOz/sZngQC2GypgaHiJ0osZi8+wqCWm0fiU8Js6d
xHCitW/iioG8KH77yyuLPj2neYN73GV4+glingW9Z2bHnEiLgWTiUKD6Gaymr4/3kr6jaTXElzhj
vIq9mCTy/rOMso6YBeW36PyCjIVbPkkYZQvR+yoAe91a3+ef3bpiiw6JerqU/O5HLc69a9T8ixjx
YJsG1Awuryy6WkWwB72aHc+g2aZORJCrZFdlzl5+1fyoRdBTi/rPK3NshEAkdoFoW2NM6v0Ikj1n
WQKw9mQ9s4O0EMDhZSGQRH4+ogjEEyUL+HQl6wXnU2ZQm5N9lmeguKFULs+g2YNOO+22lhDpS6r8
mZCbjteY6NJxV4TwkAL3q9UegLP/wMCbLxbEPK+JsU176C1Mx4snQBXOPZL+7K/potdQ08PbI2zi
S5egWddlS1GONaF/ejLcSBoftbO/p4ote2+W49WO50z9t0DxubQ5s1JmcuVdtZsF1wneVwY2lUsg
LwvLLYLHU0FXhN+b6dVxyTV0k77mSg9673AtvIYKJOnC1jKRtopbydBEvyTAwv6ZQr7JwxeubtVf
GSOxzPmurA4Q7nX2xt8T1c11wM5m7vvJ7pr6mazFJv7pPyii4ttD9DzFhCYdgs//kHnK6GDz92wZ
8slsCluQTzZ6Fj7XL83S8/WFaj9aqibaiLbHHfLDecUAM4wG/ks3D+Xh/8BWemejpp7EHoY8fVqq
L7mkIxyc0K8eCBeflz1FA9q+G5ayp2vx6whTGWtS2H7iMuLQhUisU/YvjsdX8vqFejbNcp18uECH
gSu4b6wfdM15lvUQcLf8MbiNn9pF7S7A4o2XrRSML0bH2uS0n/lD6hV3C10nyredzsaTZeUZay0O
1CkrHoNcWX/DFCg6NWtpfsoI2xMp6XYMx4a10AS3Ea/8ZdHiISInw9hUoaxGuhUFovReZm0Qwj/B
+d3D/tQId6j9iJLLd4BZTvWtMhEdm46/gkqifGluBvt1ijGYoN9y6pVrNrnW4wzp5ny5xF+F17sI
yA2DBwy86XLgm2NIw20q5NyKahRy5ZmAk+AMc5feY6AhHHokTPjFAFwQzWRCK9llkZ3KVo0uiGu1
x8WNvw20eD0ZOpLnC+N/R6GsvM77vNHK05FDzxkiUoLvqPjkvBvAZ5q6urzbzDjDv3IfgNISlbVN
InvxqPh5AiifTK+HoesypRLF2tPDrGTPaD6VzZrURT6np78n5BC+kcpEWo34obWboFP1fFgYjic9
OPjoGEZ+S9QKs28Bo8NFNzQDIG9P7ud8ouuV3vrtSs5sNTEktEHReaPuEW0w7bt2F6m1hD6G2ooe
KX2Libnzlm6Q3Ny+/9bodv288neczVGItXhdT9uO9kwMHVHCA/aI2sp7BdDNEQLLfFXj2ohlhL4B
OSqx2hR+sBJ5slv4D0KBfI95IbofQRJGMxJGwi8mmdCsIgQs9/w0c7w8041Xp0Eu7BbaSo1KCNyA
zcUXlT/uuO+cNKbS00i5b2Lbmn90+krP8KaBYlaFFx3y6f7k+gswxtzOetDfKXDEn4FHX69JJ5s1
iT8NK3XPwz2MC/PDZgtjnvmYcvbwOVj8pYebMPloQMQYgROy6dg1nJXx2DotmOeEkB6Wh9SPc0A+
rIJCrwUnmyBp6x5E1IDeqgp9jjrO0sYSakuBFGdUpopIDCLNuWq9Eei9SLwimkc7PSFpt6OmY9Zs
eZDIjhFtNj+g9zNHltcyEjQP9y7WfDV91KSABPMyfO3O8XEcMn/HluSe3YYZ2gg+MHaDHv8eylfZ
m6CG55K+LNy9knC0ta7wd3fn6yiXcNGwu7n8VlOHJjiIDUdzRaGXkuX81Gp27G97kMl3ws60XFnn
s8Lh2Mi6nC8inqqYqAnG7U4PjAq1r69eWx3fxanRx9OGgGNe5Es2ZojE3HgcpTzZOyJMTu4iAc7S
K3+iKIPxXZcH3vTm4/0G7EpPPh6g03yrBmarpaVDFpDg7vd5bqij2dBeP1PlyE48eIDzSK6LYGmT
gKkYGHdbKTXPCrLanNwrOXqeHhUI6xUp0Cg+v/It//IOOxVAEAUZ9R1VIcR5e0eEKnVKosA/97+S
Vzwyd2tSPmT6qNVAweLUgUsobmx70kAeD5fCb7WUnKBUsDM/WTwIxi2f2JUn3FFz5lwdrXRwPIF2
0VcloOAMsEhmh072DrsrzAkQuN2OHGN3fzyinj4g14qLLYrLtYCkblwwflav4TcrQFnLsdycc4Ko
xJS2IJEgieI9IiRzjiudWKiuiaKssGvTIMiO1pU0Yutqta58tUJvjptekPzHpZIVQtbIeIiA3BCX
CeCHZ7eVW3cnYSTkK/EFD3nYsU6zLWovGG4YIuiUjWjbhR/Rd7LiGSra9J5gozp2u2sgUJIAKhbi
OrLxpN9Xw0DgnjlQpiK8wX07yQWlnZqDpbqfxlMHQQBTIfmtgVozGC4EXPxzNmn4UTPF+VCEk7cN
h9aKyMQU/UxZ9D2ngU93fOs6QMR/3IMT7ssskaTafUminRvPk4GJv8IOt+Qds/XNSaXbRs+p2OCO
4vtKJOPruN2hFLdBr4l0E40Ct9qCK2hWNuX/sV3thcKifhTwnaP0uvwbp60SjT4KsPOMiQb0ajzA
+tZPUKRMoKSsGR1m7kUlGHxFJ01ZyWyAoobUkyKUoDYrK6uB/0vGZI4Hx70JMlAquGWbDWH9t4yh
IWVrXR7QEX9fLck7Yzrv4+zDL+PE/PC2gF01ExV8Eg/9FvHmcObKtVWM7X6KO6seGT7EcFq7iEmf
+7yMP9KT+QDcSZH/d6nDle+F93EcWAQ/UgRMdCK9iZBXqTF1W4U1Ey+RtgSPxb43j4hXYAPVF1ib
h9av8D5at2Mw77MEfG2SORZSR26Mr+di7/oLg0D5iFEFNbzOxfs5zc4mJ/htk1XIeTlhuO7szdby
hoQFBaynMFnBM4kaZuQXCL8cYCbaNvHQf2KysC3+NnNSBuU6O+ETttkZmO08l4EHxzR/tlxAxFOT
83PN2mCaJCfQwCvr/buvYFvPBDr4Yqb+i/7MM7rXC3w2Y1UCompTmhiAVdM5lE10c8RmTF80uQYu
TeOgES9wuxurp60wdL44twBrPdt0faiW6QgbCXZMEykMaCIQeLaR52Dt/FiM7BG1X5rZ84+Q2hBI
UpQEwZBJRUhMb5oOPSRLJd6Y8tH0V82uKClimMFVaa4E/5Q7oqbv1awDPWheRSW3/VxUjxQXtR4J
k73IMAv37GqSZ399dHCMoJhztYEYfovfHZPy9dDXfsXYI3PS6eRgkSOxPUrNhG1G5tDG3pOhvj27
y3SnhaPgavn6BCCaKUCQvvUNTVyh8Ldzs9sJtCFh2l94QIWkRy06naLcs7Vh7cpyh9iSRou0ygiu
41+7b+h5denMPbFgW0alv8wI+nCicCfJU4IS+vyfJcuYth21Z6HxMeI4cvbsOo3Kd4kaq50ifCz0
dlAH606UN+PQ23fkUD2wwMvOkc+Elr001tkPYJzgDFc3M2mwHL8Rivjb0kfh7BG9vxF+6nYe/HjN
yjoaGpNrxPly+JIFOvs8bO5+AaFOaDXZHqbSOdB1NXw9ADNM8zwF3MTZF+OGf9rPonAf8PMds8j8
Jz/EeyKawcGM3ewmQMsHXeCjB9sgnKvx3Ug0wK8IWyn6GQAfpUXrjiB7MRI34X4tv9R0Sai2TjyS
8qVIBcgFmy0g5VPdKOL8xUtgVMfiUooI890fw5zW0CbeJm2yM41zUp6PkandYy5E96gMQF4/lwU+
FxPVgP15BBdlSYjorKni/1fZfnM0xeoNe7WXT/nLh1tl5UamzOKXJPq4PEuP44aMZrUOmcXOuLtL
Xq3hHAZXnnfjQFHMDOjDwXXYaeiOsHW1YR9gFrzoNq+CM/+CeDrafjtg9IUCT9qNHYbgMlfVefDK
AZP3Z2IAC4HqMezLncxinM7wIV793sXFAfPMHkd2xfYLkr/Mw+E9yP45eYzifkFgIWuPYNd25T5z
P7IHhun4H8vqyIwTFQCv7yfw2wS9pB6bZc1wN8I0Ty80t9MnK3iWaCXgkAEZyOI+xJOPpjLhsJiS
DMWSDAynnS2nG+HeOuxvhRKZUfjhl729ha2HNezm2tpbWM9WllXO6qt2gZn5RIgIXIEjQiJ0YQGs
8i+usnZ1XDHbn8a6Ef8N3EmsgCLyZ42FasdUbS7EzNLG5Q2Di9Yv+4M7C5KZMqoejga57AiQvKz2
a1ncUmUDy5277ZAq9E4bTVS9CR/5/HZY1Swh5epPIVObsQQyIB29CfIkgktwnJS931zEk6Gtpxt0
aWKgruO8QCFh7mIki81ZXZs12ue1SK3W+EBv92tbk2dJB3qCSfnjw37PL9Ml8uybw3lB/2qzf7h/
QI8EigOMqgIpbKyco34xjmtV8ZE01tmLD+YEerhX19umH1OEWAZjDzIVrVnlvmyFpY+sqX3fs1cn
k6JuYXda8jbnl0+TuRrEBT0z0z0qk4PQPZNEL3df/PKneML9IIwcbmvZyEVO4Y+gzv3OahsNA5e+
ai5kYhudwcccNMhLwNVT5zZau5xSBIO/3Pix3HGSxmBDl2bwiHb+rrB2DIiG8zOFuAavn2yvJvy5
N/T8Mlpo+7PYS364cGzsupNaUsEmacbtgs7DdvkxH+wR5uZa+FvBJdH+bYmvITnZx5o93AOBJBFl
weOitTLTuVsFKC2ha65aiakzuXvJq+yz/X+lU0QLv6K7tXCUdmAen9HHcNWhjCN1SMXR1OIa9e2u
V+oSJgYxGOasKnp/ZZYgPQ46IhVc7U7pn5DEhyBCdvNZVD+xsYSB6EqN7f2xn3kmvFpcLWBbBKeC
VtGFKHGrzAQysn2e5WTzIvYB34tcn7bSaf2tCun/PGiNCmV9ESUODnt2H1CXmNtDFkyupVG7Ec/Y
1R5JCHsvBfN2pmijVq/TI5oQw6fNyUFu7xZho2wvsuRXUbvZBQOidSdqDzf+G8+GCSRnVQEVO8V9
oiMVek8rky5AqZFlviJ0wqg47csWtaJBxdPcTK2CLK6Wui4irbfkbHLBRD/G1xCgyzFEy8gT2yIH
6or2bZNkkPfYE5/iLms2BqLf22hFEv5eVy6Tk2tqiX5cjp4RQtcTEp8Ot8upsltJ8HPvdtIwNaMl
/sUtplPRZrJ6BcgvJtv31iQHcyMsGNqhZdOxZ84TMGvE/IRCTISva4fS1YtcQOCC/LL+nRK+g7z/
FwMayELU6xOf61LqunsNaewMtcYpTOAVcochQxhiulgN/1QWQ9gQ3TsUuW2I9INuy3dgpRGSNIx/
Fq8p2MJoklRF9PU7kKSma8UE16NpGekU7lXy4O1g5rpuDLz3GBgN2dhMGX8bhzlTzRynqEy++od+
zHuGS0Izy4+AjAuaOzpszjg9GlLxkjK16TPsb7fq1jn3LmYf2i3C/Qm3o2r7yL1a7gzsQ5W9Nc3b
x6Vn3iq3xkHflmGV3Y4z0zTVeqebCDaRrXpqQO7mDP+PyoRdDQFGBxv36opPO3tulPNVuCL5BYAH
2lFQGWjSyVhj/Mj/M7lqQrw8yMiIGyQZAyEP4DUo6dJmgBqIRrZZ8Dc/N+7lxFxV3hdqSwzV6iWR
HzGT7U9Tgjwni5cdAIvh0r8vqFSTEtbOidmAhETX01Y37Cl9j39hkNdraH7ix7Ph5npkC+Hi9LZk
n7ezlUmZuchVUm7//oSZC8lcW6nrpIZxQgbdU4ujxvGK0uq7i75mjwVievFNS0BDkBOxka+tAt5V
4Z3P6MZvZ78k8tQqD9bC2fbTgerVUtf1tFdsJGqV+0Gp5ce8dCwKn94fJ1ehCgE0CBZoK9m6JGYO
P9qkg/ILMbqSLzYvPqi7dttp/2i329h2seQSbi1PSZt779vne6KdoWROezXz9AZqnr8GDmqMPuwc
U1AQZdJ2fkZduUJYTpQD/IEgtegOIFREjPX4hNX1/yrYwrYfFCQ8syhXs2ObokeA2Q1/eYJUOX+W
dVhQtBQwvkpp20ZWLo7WLQQhmLTCxZQNQipEJsYnP3HEFMK78OPEpEn+zPMhN/sk6gGsevWyK8Pe
q7BFlPLykpOWfZUSCQdxdMfoOALKKFAzXooBrXsF5O3qa/fmaegBdunsLyOQS807A+mtJvOe6HH1
OWYz1mc98gUWo6McQQektlBVAgSE5ZWYmfMINGYPXoqRbv2hGD3CfBT9CXO4sGQXNE8X3i4C6V8O
GEx6VIGj3Q4XYWkjWwh3UGpF2wknyyG49Buj8wBvHxcoSxgZh6U411RhW73PGlsHkI+Ro6pJVGsl
bBddH23ihzyj1ZxVrnHXdKg5vcVPcbb6wLbv6JWdvoe+WqGuFTKcuD4pzKq7A/UvpKdi9Oe3Ww/s
By45H6xE58sdt1MWULRvYhCK7ig107b1bX07aQ0pcDtdzscsvC+y9m7NIGK2XC+ql9IQqOPXkoUq
9N7OtOfBz7KCZeFOxAQ39KBhWZBYVxUhumXytKmg3TStxXCuLBhCHg2L4ydvBjUIaGFisAn6pgsW
aUeZgg8XPyePBRz4VMGwLkqQuJYpdmDpDExV1zrtbf8rqdVIwXw2aKqtsSl4ZxeXyJI1pPdvKM6w
msTWUGcU42LnjAOf0PM8VmP4FWBLYWtJFVZpB35NSBGMXJDHJuku4Ju53c1y5CN6w8V29C8pPjvU
rL7eBySz/yDggM2+fI1y48JIDfpZuYNWE05u0ZP73hvimaymAgr/+xOYE3yNiL7EReTz6eWO50zc
wu7RkkJbeeWdTyPL65kX1wyHf1YPalGu4arMilSQI652uYTHezd6HhU59kjG6CKrgVUEGOqb8Mw7
5UMod9m1D8eK4SRwqwpy3/uapH4UWttmTMLOdiMxRIsTs6nBPCOP/iXsZwSqU/B2aVlCFj43h5/c
59jCAik3cpw369jhYihKqcyBXWmU7yK+uDW9njh83EwuX1FD4M2FMRrFV+5RCO8nP+L5Z4Hb7S+d
0CFqtwjd7fI9rE9+GnHUqfEvFuP4XqdBwWln57E9ToVZTCk6cil4vm9rbxwKD+PmrPM8AdW3RoO5
B1H4qEbEWg5vf2Hx+q47gODisoIcyh0Zv+l5fWep7JhczT4500bbCRsny5YOtHs0b02iyV3eAjuP
/5b9L412wG3xIGIMiyNK7OIo0EZGgp0rBxo1vyrZZketqXbC/GQMh5Qp+GCfeWaJUDx/vaWJVBjo
aDMtV8Zv7yeD8GiO9t47RmWQCutWmovf0+HHFBducPkLMEC9CcXkWabHuSB8lbJRMTlvU7pgtf8e
rIllA+o8UWW60pGm17WMl/D0uxeJLa2iJQO3kyOa218xfCI+nDdpK7Zu88lgCalkl2C3FtgdcH0z
XqAhKa9s88OCZ+zBUYQ9GcJchaHxXx0lkMulyWPPrfODJI5RVswQiAtUpPoo8zPzgC4+sStwqwcV
WRK8JQQ41z2O7vfz/qFNMlZDfYjGyPC3Tbmy4pE1XM4iWOvqm2iGUMXZXZQEAkYGt/jPo6sreQSm
WehxcoAXDReurwzWWmfGK05p+QsWKoeWpmBUnbZKJqVIfnuhWvNBp1+oGF2prx9euEzOcjrMnPOG
hNhN8jXSrJI3C63DycNbjhV1KjPhFHIkR8N/TLeg3M3O/D3NocVAfIe8SNBnXbMwmrErihzRHsrY
ppJAtmizVpKGbcL8ITXd75igLOZgfcHwTiGrszQsws8oo/OISObGje355XZXtkvWhki5pZnkW0cW
3ZXQD/SlydzAXGRsekt7vvrXbHpWNNHcd2rWbUL65cHcKo1GADXkPVGebbavpB+f/WeKtcQUWtDf
iBZKzr1QE3TT6CSuzeG/fvvrAmWFxPf00D9vEC+tgQ4L5Y7hSfWkCmBadtKPYOEdKQj5lmyote52
0S/DClKYt27gYLuzKrlfX6PxoQ9xayMLVNiBrF7wjCHyFTYQPZ2owb058+Fj47WPx8L85Cz/FU3y
q/n/7rPvwF73s2s3qJ2FX+nS6ra/sJvWFdT8BNiVXSBU1IskjVU+JmWON4ojNOrnQDMvRLEDdQ3Z
z8H4O4+kT1G2g4knV/NRXQFCVI5BvHzqDvHZUGp5U5wxmHgNf+p2zKKsz442d0SozcrK/RAw+dMO
9i5GN2Hz+3ASaMLx2eeaLNHcppon991HWeHBqmqkWnw9hHb1ZL4yUN5qnxmVDt1VMkymjYunCQm9
NLpZ9QItgA6FlK9mIziPyiQF2NbnIwg4DEY6sgfljlzI9fcdfsBaanomhNJK3bDpHdsm88SY5X2i
QLmM89q+3CzJiBzT3QC4tQjXVcszQvZd2/tM/g501LbsyI3jN14856zv12IW4cSh8Xyg9WLmsbTB
efTqjX30Pm9kEu2gho9nT+hJzWGqD/nkdTlgKwvakpW6zIh6heY7SppYF1CH9RdqVOGYHG9NaM0T
3SK7h+mvJVJ3tExqoBbBo+iq0UvSOdrp7UYhcF9yKKqGv7hj0I7e6iD1HFucGpXwMeDqjvg1ZjwI
P1xJ/0LX6N2cps9wztaR5FPEirvI9lem+5sammzHhQCh+JRhFxD1ZkOI2LVylWnsVaXTXe472DJV
J77Qd71EDA1odd7OvQ5Vev8Ztbg1sOJ89rfofoEH+uzCIwA6Pf0pmVIEB0SRkHvIiNLtRZMdCR5J
eIDXlpafswh7M4lOXHhYKKiLF4XD3b9Utq40CpiH4h4mNiImPkPvo2dYC5rZZDiuG7iuB8Kuhg4r
eT20rtU0XVF+Bd+YhnjZ+3DUtbr10mGNrZ2HByI+fkHToLYz6Z3R/NnYczOgZYee9OmD3sR5rWFW
MuABPYDocER7dwBHRUb0hqmae9SE4Ffx3FAPgz+RmU1zqBSy5lgiqI4Y5ykFNyeVLoWoZspELYVS
QvVZI7sip4ohJcpNyyGohuVidf7oipqSG4x8AAq8P9HIMXQ87qQ3Pb/YVOL+P3oxa7JFlc7b1bkh
oYj94LW0l88ia9Vb9obCeyOLL9hOyX6/uUUeaTphpW9pWkxLSSWsWvCz63B6igvIhE4g1v03G0m0
g22xVEdZVMCLMcsauNYdBQL33dsZRa93IpBxApb9ZEm1pvDKVkwR4/qq5X8S5fiYPzhJ27dG0QP7
ykuP24742zZtN2OiCk7JhTCA0juFx699HWLJALlxoyZfvbWcDGpV0mUNQZ8fx018w68E2dQi6AYB
3x4yMprk10kf3L9X0/a3YWitkeXJmO25FFt7sT+34ef84r1hoHZoeZmyO+8acdi/7xq/jMTKTuOd
U1++IFgMkG+ex8D7/jQIjZaMdC9FCJsF9YeEliLOgPCQ8okHQV/ApZCd43haYU1Tz9gb1Cu1iaen
8175Jqsh7XVxsx13RRorKv0RAAbqFVdttEN//qp7D1GuohRs/+2ql0YDKIZd+2dIivaaWONafJaz
Y3HxVBXNG1++j1ymt1wHgRJKHBfrfNVRzSfx86Wxmh4DFdAN5eDUOqqHAnzEYSzM78qILBkWIjVj
yEZF9yctWDXMVfQ0zmQGzSu8fK5vF+UsQUxwx9KBj8xPFPYyCKnNlHcvBPiRxGrxoBdp47NxyD1/
IKcVX1xkzqTQC3TPnX4iJy/xjhYJ2CEhJbFO6Pa1JwSm8IdHHSlLT0rIaSPviAFUQ+k5LNyr+j5E
DBRs5u//IYsnloVVYGoy9UnTaUDnbdan/0lObxIaO6IlFhQADkmkuIBtQ24VrRcKSR0lbj7VKOuY
LLvQ8+6fWqTg+m13mjZ372hanGoC+65Yx3q1tOu/EgD53/qWGsp9X6E4HIUrEawa8E6WvIQYrYb9
QmtFDet+5v9uepPS5Qy5MTTCvHOZGXTiuXhr9bKsWRaC+2BKBOaSyXdjVX3tThj4MEUxYSgaIdX2
abIgsT1gTyBa9gK7aez+hCOdAbqur/6kMA73aEm5knAIGv/Mm3NiXmwZ3if3lDjVgo6LGhpArT1X
uZX4R/Y/SjtzXpwfwNsCKVuMTUfBmMud4w3p586fKzTdgTQHN1B9A2OxqCDpUW4LZdWSBu3lhwzM
bclPW1SAYq7Cw10QNnE7dlCz7C2h6H3J6ju7CRBRcCN1X3JYPCaJmhkgltXRNsQv1BF2du+KNm/W
Vd1SPJslemAN0VJoVJuwS1Sv/ddZRf1FreIgo6nQkSTkLKUPWfPV84mwmjrWz5RD3y+fc928XcnL
ba6rKvn6/yo+yzfnM1VwjjAnWXPprkKT8rSm0dDseukJj/WushMDE3fZuWuQ1Iy+Ifcqfp9VuKyI
sGqWGmzKvUVOhKmys73cHKlkvtr9WIFTmNo2IT1zIDTDIZNlQrkNTW0zxrJtiLaTiGXlBv3RYHzD
mRds39+p4mDldw4s9x4hS+3Ode/41yaV9JU10hObd/YWT/K1nZqI6XQh64vshCABaopiO5IoclLB
n8JVQRYO/uo5TN/5z7BTUPSZGglNlWt/q+LbRFY2OfbVXCoZebCXNyzTejDrgtFxIJBEgXZ9W6mc
A2QYJ7JSn+JMZoSebSPIvRW9ENMSJXrtjegw4E9KgzoXLP0qmHX5lNwOxNxXILhrS69W+Kmtq8CP
YUJ7Wne+kYYnR26MKL8kmNOW8835Ob6NijkqiTi3nOsYoU3Zikf89PC/njtbYmcK5qMSDdMXqDjD
qQyoJJl5/Tohj/MWkdOzmtsvLLPJ4KBw9rVclS9LYpWLMfX7KlbCo9kdweaBqmCzwCap4dMqrgIY
MbU6+YWe3kEkFWdCUsB7OYpgol81zyNpGypwPt3y7MkZPnrvovE3ua+Owo/XpnAwogkvkVCL+QpZ
3k9+jwMHjNH18TyqeFcFnv1bpCa3qhvMVbgABR/VGTD0dedUvV1TsFRtD5fSIo9GRGUH+4dE75sU
6q/OxncdXs48I0eYmdRVbvtcgotZYu7SlW9jcPsfiIpg81iRqxm1b7zgGDkf60+CTfnb2d1RZKmc
tpCjXYmVe4oKvPsI+TinZQ2K/pU/YeL6U9OZ05ygVNuYaRFTnGBSBYoFqzzLg6GTV7D8g50fHG6D
YBlHXSClktAF0gzpAVvpLNfZsHidlBGnza6kEDguSvD7AUidicNDjmFyKVAA6pEHRd4rWypLHR+2
6PYY1PDWRUVJ5MAD1ooHKjWwcwCqFuhFDlm3b0xllBf6dhz/AhBbLxckTxokDc5GkSpFFUsY884q
vu69C48ssrCxsVQOSycHtgiojtO4NhItZVvMXeEadORGu4R66/GUeQ8/yO4fP6EMQ5K0r5g4PQdU
gZa4ZSOvSwcmjaBewjNUwqWf0XNKUVpOkETslHK4h9VPoKeUPFsL7juzv3tybpNYfN2bAkrlpWBa
9Z0BWMk7SVhpewlC8P9qIVsraEZJw7tWC3ETu8JEgftS6kBTPkDNSNLhM9oq+jDyJmS+4bPZhm+6
mycRrmYomULVXbm8vn7TOIzqRmkH4URO4Dh8JcwvonI/v2R4y7QpaN1mNjd7XpUd6eH65UveTKxx
KWVXNWvGIqVJl7/8sdxmEY1QyEgPsVvCtRsl5virHsSFyhahgI0V8XOsVS4M6UZxbYPXPtYLftMi
EYdESSpJLC9rfcOKiPkVkiBdf/dGkddFRe6Ryr0hhY4cvYPG01bBqZy4yOyVTfzO2J5jvi2wtCEm
4FMe/OrR1hvMu40Mc57O6Ue0J0r1rxh77WK5ePSBlQ4KH14xXgjWL3N0RQ2UAAkrP3HYPaHY6Pyv
hwCxMHbmAKVQxHE0UoCDC/P02E4fHvBVcF99u70SU1xxCdnNA1qBB6iUZRftmsvgPX8iOzeYDFvy
48oh+SXGt23jKAmSVksaQTbK1fA1euYyqqeS5uTB0OZZf1qYCPFi1MmI9tlBZrVVOrT+X8CG5j9m
6PAfzv5zRNXv71+BY4QGcva1RrpOGPN7OX2vwHCIZpwwrKqtgeeYYibt3RK5tW1MdyT+21PlD/8A
RiQDFvetPJg5Y5tbPQAIBB0Q6I6K0aIBT3vMiZdvR3rXgt/k8f53WpuIGJYL2Y3aFb9/f8v5uHDM
sPNjuMsYLJ+LW7ITQwlWk3Si2HD0DVecuqhEZ8mkdnD1/h9tJGWjYIEp2hzghlRUsBv9hYG71VNP
7nBlOzNle+CVkt4F9qu0bIHu5MczT/UpyLBlZIEC0UxoCYBYdCnrjdb7GyLTv72zS3Ocbt1aupY1
eu8AGQHAHitMJi08mSFbMZw/UZNiSeTshz4nvg0/rgmK7m7+28V7/HG2l4uuIU7qsq+Z3RoeW8DG
QPX2WnEN7oYUU4lRDsfPYBhlOxkm4sEFlJ3Q1HnkSXIMAWRn/67V97UMlQ25bDSQwepLwv/o1gEj
LOwcNSMxiQ9r8FhhXDva59rtbT1JUICrdgH+wyyWT5yUn+WtfEPfNsejw6mvDwGqxRnfes5Kl2Zv
AKNjb4kEZC4NSQR4Tv7tXEfT0cjrC0BeMTDyZUhRHDIS4+2HcxVhRgsC+znb/pQBF4MPGfvPd1ZV
pqtzICnaNqjH8tTQo3x171L5jyl1bChnnX4azVJHraGyEw1uyTYKfu4UxkG16OV8q28JTh4Xn8I3
7VSWCMQ0mLM09UQO1FihIVqQZiWAgizHWQN3k6UnRyjrCYZdgCtVyfR6D1sLt6MfHCX8TiRSIdYT
W/mTTjleVGaPm7c0Aa5Ws1nuYmXKzze/SiW5qH/MgvA97zjUoZtl3c5GecE1OCIg5XJqpam5p3CE
NEXmLVgCdrZRojpq+p5DExJrWEnMawm6hGDY9zSKAuPj+Kuq6JWPeU517XVfREKrj3xTTCdoAp5k
OYZGA2JFfzdqcT8B17PMOrMfpWGK4KabZPfIlSxYf+jCpoatvzxf0JrVhSmtu9xkOlbT4aos+KEn
p2Oj9Mh8dFbivfmcB+ilqsvU3vCozy2tusyuKIEpMVb4560GGzOJGv10H/1S91EgfXJFKqg5JCoD
aXW/XjLtVXa6lLCTOzd11CWLPVYrX861uZKWwpnrlWxw87GdWvdrzuOWWPqdAYms+VXDk/Y820Go
bDxS6D0zVGDiDWM22apbGTIbi1LREnD8rWRVxczfiiE8xmzGI+RFIIu2Zo45J2l5thMuSPFYyf50
buHqhlrzf0sgI4HXt2tUssO1+5SDuHT7bGCnnTJu+fiiom7BPAL5HeJ6jXgdtamxA6axzqv8Yl7C
FGxFvPoRVcbS/kp0iyRL/JaJV1JZCECTn/cFcRGUAimKr4hlkZ0pafZ6d+8WuSIgl+pBRDNWoRUO
7JCGDiHzKQW2BeD7OsufBhJqFlM3knZu3imQeXfEwyJ5NkDs7WN4KaAiAbWBUW51OS9Xdjh6gvUA
lNX6hR4sYu+vcedvqfIyn+O2AivnV/UM9wB8KbCtP/Y3/mWbR3P4JpcId5ZgtmUTGl4wpjpLeYKw
00JCaUAgcFYT+tHUOaek9CvjGQjyr8qKPgis5+IAPx0wtGiWFB3nARVQStzwh69OrONN8bdFEWfd
5ph1eoaqNIFwpF7b6GT+12OQhMbn+DAhWJLcYsZQ2Sg853WgmFUYReBJkTDHo9DHCxmvFJh7B3kd
fD3DssmAsczkbphfEXPD0/uECMq3t2YgYiUrd/cK83buc3ciBYfD5iBXO/9dYN2zjeIw8tSxzH+/
hxhBChp7k3AeCCS9E5zMZSPyYBgmftEzH/0e5t7o3eV3wHMBmcbzimohbZKMbhNuujRzOMD+3DtB
sBTSAVBEvYOMxbFJTZNu1o/kHrwatiz53zQ9/4b4+yDt18qgnn/zmDagSy6FzGvGd/xSc0fvMQos
5Q9bzTgFWWEDOOUwh6UmBulp/PYWwohi1uxWtG/VjccXKYvTfRE4cx6whTxF6hwmXrDNplCbBGlO
3DBPXMV3aFmASmbR+KQX7lT4BGBKMo3CfIyPRrNa70W6ToWDYW92BgX+MSGOiifoYRIn7yE6zp9F
imCcpZWHL1apC4B6nF9rqciCqqn/rpTHG3vMKm/EwEsF4kH+NdDwK1APlp3dOzeAfkpSxrAQIo3e
gjAa29YrtS8MN/uSRIuEee8j/c4d35HqSOCawLk8azAIJdE72gf4U7YVEpYF+5slL2fIRRZMOd4c
i4seIvvDcGRTo8adRXVPxdTy939QmWfbrLuweZd/BtT+NohupmgMCErXUhxh/BG4oDtOZC0EbYTY
af49Ymc/pd9kuvuEz/gdNKRK7D4EIKUo8nqHe9YP+uzk1NlFF7Kh3gEZgjCMA+LRpY3r7jQqrrD4
kleR06DNh9avb0U1cp4JPNf3kKz0wKXqb90hz9JyDF30dYYOAPVwflH98bb2SHav3ACLwhiDY+jQ
wE3UVWe3F0PFm8LdHu/T3jqGj5yqOmE3lzO0B+kYjVU3E+SJ9xN7Uy89oVeJA8f+gPtZg3vVL0pj
b9/CAWgEQyX4eVI99dq/VX1ZDtf/85ZwZJ/UItaQ2ylQKR0abk/SCJATzD9mBNg0GKRqiUta/SgE
iXyuhO2A8gSbLXliHkiPnA4eGQMtRL/MCS14qS/+bP2WZIWOOcKrFumiaFEwIz9hu9SVsoTz5HoD
8JCV9pgpMLcr9sM1yv/KNwYicMAqjVvaeqcbdvTih3hvqfj6tVZBkW7uPRwYD+IC6AIc4W5xzNRP
RkBCzEsAtjbitzUccHWTYTWbxmKXs5q0taVD8da6sqvwqf+KysKs0fMHu/ABO3osanSTMvThhnU1
iHkwUq0nk7jhshDy2ULWCu46mM5Bu9MRXU+i7bgVOoNEdScTVaKmoJm1U392T9GzZp2T5S0qGlim
5O1kEGFUD9YzUHyD9wm7J2Pbg1z+PGlZT8+fuvDik5aJ3Tk8KAzInIHYY6IdMrF5It1bk7yWY4Fp
+rx6oSIiB3EbH/2TAlHauLcAL7Cak6HPVPRfFHkcwwwUrzll9lDohPJOBYICwg429zAB2kUXQO+0
X+RzRHTb4mC/iCsseO8oPU17JWEWP0LioEcHMROA+/KyS03xU+4p9+a3GCjO3UX0cij3tH1TOPfP
pL31zy4cR7reF+qjl0dPmwXlBoErIDVnmKzbaXs0ZNdU+guSR84vLQvBt8E1BIAs0vqoD2lfftAg
KwPCYnE+fPBlYey+KbYzmBfKh4gmS9yuUz+G9pdI9U5/r0zwYilbLSc+9F2Ro7ErIkHmm8/7t3ez
Q+fP1zzS+0XdBDSwj+D7cfB4fV1t89zPYgkrkQVWsdWa+UEJHA/JTn0e8ibVwueZqZePDW5zqNAK
bKcaubQCZb4CqGh4K7p1JvaSMYGoygoAPxJDkBClbrFjX5S3tfM6dLIGSe6iIJ2jhSy7IKYpQ2Bp
VN4emPzwXVJJtIsAonut/NOMT+AX1M23fxygCDi0puz7qN45JCTN5ZI80u/YCzXV7Ns2NdkohyBF
AFH9UNV4cgry2SAEiL1VSWV0D2EC+tlRt1wMmbFPvAnqO6cCJnHSmNS8O7sFINe+0vyMFUF231lh
n5lcamJqhg47tK+UYA1VATcKuZLDywfDI64UTuzBUh1DHMk7Y4QTfCwUdpQWuFkqx+5aMSOzgDvQ
X9uvAZhmAtIwUfS5njZuiYHpVi6jp6dKfA3B4FudLgI8Lin0h6iJKCM5bY0V7sEYnn3ijRQEfXLU
8pR5/Orf5lE0WaEgbYDlgsothsN/utRN49mh1ZWBufRVb9JOo1vbzrUx5vGaKtZuuhwrUALk6P8S
1JCXbzbtIPLtM2kUTFu1dho79RrLAZsJ4Y3cQhrpbJA3aZfRUwuZxloWe+LH1IVrzqUlbK2cqSHY
LN8WprWsh08Bw3tIryjlCpr95Qc2FmXgybWNC+VLNWFCocF+EHVoymiV/Xp0Oqsi6wQs/PSscH+0
7x2x/l/nUDJPgkSFb626AWaIGyRXua4cx9TByXrDGzUnTQQskFmEP/Z365ZXm4le
`pragma protect end_protected
