// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 15.1.0 Build 185 10/21/2015 SJ Lite Edition"

// DATE "06/24/2017 09:05:46"

// 
// Device: Altera 5CSEMA5F31C6 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module sine (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	clk,
	clken,
	phi_inc_i,
	freq_mod_i,
	phase_mod_i,
	fsin_o,
	out_valid,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	clk;
input 	clken;
input 	[31:0] phi_inc_i;
input 	[31:0] freq_mod_i;
input 	[15:0] phase_mod_i;
output 	[23:0] fsin_o;
output 	out_valid;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \nco_ii_0|ux122|data_out[0]~q ;
wire \nco_ii_0|ux122|data_out[1]~q ;
wire \nco_ii_0|ux122|data_out[2]~q ;
wire \nco_ii_0|ux122|data_out[3]~q ;
wire \nco_ii_0|ux122|data_out[4]~q ;
wire \nco_ii_0|ux122|data_out[5]~q ;
wire \nco_ii_0|ux122|data_out[6]~q ;
wire \nco_ii_0|ux122|data_out[7]~q ;
wire \nco_ii_0|ux122|data_out[8]~q ;
wire \nco_ii_0|ux122|data_out[9]~q ;
wire \nco_ii_0|ux122|data_out[10]~q ;
wire \nco_ii_0|ux122|data_out[11]~q ;
wire \nco_ii_0|ux122|data_out[12]~q ;
wire \nco_ii_0|ux122|data_out[13]~q ;
wire \nco_ii_0|ux122|data_out[14]~q ;
wire \nco_ii_0|ux122|data_out[15]~q ;
wire \nco_ii_0|ux122|data_out[16]~q ;
wire \nco_ii_0|ux122|data_out[17]~q ;
wire \nco_ii_0|ux122|data_out[18]~q ;
wire \nco_ii_0|ux122|data_out[19]~q ;
wire \nco_ii_0|ux122|data_out[20]~q ;
wire \nco_ii_0|ux122|data_out[21]~q ;
wire \nco_ii_0|ux122|data_out[22]~q ;
wire \nco_ii_0|ux122|data_out[23]~q ;
wire \nco_ii_0|ux710isdr|data_ready~q ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \clk~input_o ;
wire \reset_n~input_o ;
wire \clken~input_o ;
wire \phase_mod_i[0]~input_o ;
wire \phase_mod_i[1]~input_o ;
wire \phase_mod_i[2]~input_o ;
wire \phase_mod_i[3]~input_o ;
wire \phase_mod_i[4]~input_o ;
wire \phase_mod_i[5]~input_o ;
wire \phase_mod_i[6]~input_o ;
wire \phase_mod_i[7]~input_o ;
wire \phase_mod_i[8]~input_o ;
wire \phase_mod_i[9]~input_o ;
wire \phase_mod_i[10]~input_o ;
wire \phase_mod_i[11]~input_o ;
wire \phase_mod_i[12]~input_o ;
wire \phase_mod_i[15]~input_o ;
wire \phase_mod_i[13]~input_o ;
wire \phase_mod_i[14]~input_o ;
wire \freq_mod_i[16]~input_o ;
wire \phi_inc_i[16]~input_o ;
wire \freq_mod_i[17]~input_o ;
wire \phi_inc_i[17]~input_o ;
wire \freq_mod_i[18]~input_o ;
wire \phi_inc_i[18]~input_o ;
wire \freq_mod_i[19]~input_o ;
wire \phi_inc_i[19]~input_o ;
wire \freq_mod_i[20]~input_o ;
wire \phi_inc_i[20]~input_o ;
wire \freq_mod_i[21]~input_o ;
wire \phi_inc_i[21]~input_o ;
wire \freq_mod_i[22]~input_o ;
wire \phi_inc_i[22]~input_o ;
wire \freq_mod_i[23]~input_o ;
wire \phi_inc_i[23]~input_o ;
wire \freq_mod_i[24]~input_o ;
wire \phi_inc_i[24]~input_o ;
wire \freq_mod_i[25]~input_o ;
wire \phi_inc_i[25]~input_o ;
wire \freq_mod_i[26]~input_o ;
wire \phi_inc_i[26]~input_o ;
wire \freq_mod_i[27]~input_o ;
wire \phi_inc_i[27]~input_o ;
wire \freq_mod_i[28]~input_o ;
wire \phi_inc_i[28]~input_o ;
wire \freq_mod_i[31]~input_o ;
wire \phi_inc_i[31]~input_o ;
wire \freq_mod_i[15]~input_o ;
wire \phi_inc_i[15]~input_o ;
wire \freq_mod_i[29]~input_o ;
wire \phi_inc_i[29]~input_o ;
wire \freq_mod_i[30]~input_o ;
wire \phi_inc_i[30]~input_o ;
wire \freq_mod_i[14]~input_o ;
wire \phi_inc_i[14]~input_o ;
wire \freq_mod_i[13]~input_o ;
wire \phi_inc_i[13]~input_o ;
wire \freq_mod_i[12]~input_o ;
wire \phi_inc_i[12]~input_o ;
wire \freq_mod_i[11]~input_o ;
wire \phi_inc_i[11]~input_o ;
wire \freq_mod_i[10]~input_o ;
wire \phi_inc_i[10]~input_o ;
wire \freq_mod_i[9]~input_o ;
wire \phi_inc_i[9]~input_o ;
wire \freq_mod_i[8]~input_o ;
wire \phi_inc_i[8]~input_o ;
wire \freq_mod_i[7]~input_o ;
wire \phi_inc_i[7]~input_o ;
wire \freq_mod_i[6]~input_o ;
wire \phi_inc_i[6]~input_o ;
wire \freq_mod_i[5]~input_o ;
wire \phi_inc_i[5]~input_o ;
wire \freq_mod_i[4]~input_o ;
wire \phi_inc_i[4]~input_o ;
wire \freq_mod_i[3]~input_o ;
wire \phi_inc_i[3]~input_o ;
wire \freq_mod_i[2]~input_o ;
wire \phi_inc_i[2]~input_o ;
wire \freq_mod_i[1]~input_o ;
wire \phi_inc_i[1]~input_o ;
wire \freq_mod_i[0]~input_o ;
wire \phi_inc_i[0]~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TDIUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \~QIC_CREATED_GND~I_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ;
wire \nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|Equal2~2_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ;
wire \nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ;
wire \nabboc|pzdyqx_impl_inst|AMGP4450~q ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0_combout ;
wire \nabboc|pzdyqx_impl_inst|comb~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ;
wire \nabboc|pzdyqx_impl_inst|sdr~combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ;
wire \nabboc|pzdyqx_impl_inst|dr_scan~combout ;
wire \nabboc|pzdyqx_impl_inst|KNOR6738~q ;
wire \nabboc|pzdyqx_impl_inst|tdo~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;


sine_sine_nco_ii_0 nco_ii_0(
	.data_out_0(\nco_ii_0|ux122|data_out[0]~q ),
	.data_out_1(\nco_ii_0|ux122|data_out[1]~q ),
	.data_out_2(\nco_ii_0|ux122|data_out[2]~q ),
	.data_out_3(\nco_ii_0|ux122|data_out[3]~q ),
	.data_out_4(\nco_ii_0|ux122|data_out[4]~q ),
	.data_out_5(\nco_ii_0|ux122|data_out[5]~q ),
	.data_out_6(\nco_ii_0|ux122|data_out[6]~q ),
	.data_out_7(\nco_ii_0|ux122|data_out[7]~q ),
	.data_out_8(\nco_ii_0|ux122|data_out[8]~q ),
	.data_out_9(\nco_ii_0|ux122|data_out[9]~q ),
	.data_out_10(\nco_ii_0|ux122|data_out[10]~q ),
	.data_out_11(\nco_ii_0|ux122|data_out[11]~q ),
	.data_out_12(\nco_ii_0|ux122|data_out[12]~q ),
	.data_out_13(\nco_ii_0|ux122|data_out[13]~q ),
	.data_out_14(\nco_ii_0|ux122|data_out[14]~q ),
	.data_out_15(\nco_ii_0|ux122|data_out[15]~q ),
	.data_out_16(\nco_ii_0|ux122|data_out[16]~q ),
	.data_out_17(\nco_ii_0|ux122|data_out[17]~q ),
	.data_out_18(\nco_ii_0|ux122|data_out[18]~q ),
	.data_out_19(\nco_ii_0|ux122|data_out[19]~q ),
	.data_out_20(\nco_ii_0|ux122|data_out[20]~q ),
	.data_out_21(\nco_ii_0|ux122|data_out[21]~q ),
	.data_out_22(\nco_ii_0|ux122|data_out[22]~q ),
	.data_out_23(\nco_ii_0|ux122|data_out[23]~q ),
	.data_ready(\nco_ii_0|ux710isdr|data_ready~q ),
	.NJQG9082(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.clk(\clk~input_o ),
	.reset_n(\reset_n~input_o ),
	.clken(\clken~input_o ),
	.phase_mod_i_0(\phase_mod_i[0]~input_o ),
	.phase_mod_i_1(\phase_mod_i[1]~input_o ),
	.phase_mod_i_2(\phase_mod_i[2]~input_o ),
	.phase_mod_i_3(\phase_mod_i[3]~input_o ),
	.phase_mod_i_4(\phase_mod_i[4]~input_o ),
	.phase_mod_i_5(\phase_mod_i[5]~input_o ),
	.phase_mod_i_6(\phase_mod_i[6]~input_o ),
	.phase_mod_i_7(\phase_mod_i[7]~input_o ),
	.phase_mod_i_8(\phase_mod_i[8]~input_o ),
	.phase_mod_i_9(\phase_mod_i[9]~input_o ),
	.phase_mod_i_10(\phase_mod_i[10]~input_o ),
	.phase_mod_i_11(\phase_mod_i[11]~input_o ),
	.phase_mod_i_12(\phase_mod_i[12]~input_o ),
	.phase_mod_i_15(\phase_mod_i[15]~input_o ),
	.phase_mod_i_13(\phase_mod_i[13]~input_o ),
	.phase_mod_i_14(\phase_mod_i[14]~input_o ),
	.freq_mod_i_16(\freq_mod_i[16]~input_o ),
	.phi_inc_i_16(\phi_inc_i[16]~input_o ),
	.freq_mod_i_17(\freq_mod_i[17]~input_o ),
	.phi_inc_i_17(\phi_inc_i[17]~input_o ),
	.freq_mod_i_18(\freq_mod_i[18]~input_o ),
	.phi_inc_i_18(\phi_inc_i[18]~input_o ),
	.freq_mod_i_19(\freq_mod_i[19]~input_o ),
	.phi_inc_i_19(\phi_inc_i[19]~input_o ),
	.freq_mod_i_20(\freq_mod_i[20]~input_o ),
	.phi_inc_i_20(\phi_inc_i[20]~input_o ),
	.freq_mod_i_21(\freq_mod_i[21]~input_o ),
	.phi_inc_i_21(\phi_inc_i[21]~input_o ),
	.freq_mod_i_22(\freq_mod_i[22]~input_o ),
	.phi_inc_i_22(\phi_inc_i[22]~input_o ),
	.freq_mod_i_23(\freq_mod_i[23]~input_o ),
	.phi_inc_i_23(\phi_inc_i[23]~input_o ),
	.freq_mod_i_24(\freq_mod_i[24]~input_o ),
	.phi_inc_i_24(\phi_inc_i[24]~input_o ),
	.freq_mod_i_25(\freq_mod_i[25]~input_o ),
	.phi_inc_i_25(\phi_inc_i[25]~input_o ),
	.freq_mod_i_26(\freq_mod_i[26]~input_o ),
	.phi_inc_i_26(\phi_inc_i[26]~input_o ),
	.freq_mod_i_27(\freq_mod_i[27]~input_o ),
	.phi_inc_i_27(\phi_inc_i[27]~input_o ),
	.freq_mod_i_28(\freq_mod_i[28]~input_o ),
	.phi_inc_i_28(\phi_inc_i[28]~input_o ),
	.freq_mod_i_31(\freq_mod_i[31]~input_o ),
	.phi_inc_i_31(\phi_inc_i[31]~input_o ),
	.freq_mod_i_15(\freq_mod_i[15]~input_o ),
	.phi_inc_i_15(\phi_inc_i[15]~input_o ),
	.freq_mod_i_29(\freq_mod_i[29]~input_o ),
	.phi_inc_i_29(\phi_inc_i[29]~input_o ),
	.freq_mod_i_30(\freq_mod_i[30]~input_o ),
	.phi_inc_i_30(\phi_inc_i[30]~input_o ),
	.freq_mod_i_14(\freq_mod_i[14]~input_o ),
	.phi_inc_i_14(\phi_inc_i[14]~input_o ),
	.freq_mod_i_13(\freq_mod_i[13]~input_o ),
	.phi_inc_i_13(\phi_inc_i[13]~input_o ),
	.freq_mod_i_12(\freq_mod_i[12]~input_o ),
	.phi_inc_i_12(\phi_inc_i[12]~input_o ),
	.freq_mod_i_11(\freq_mod_i[11]~input_o ),
	.phi_inc_i_11(\phi_inc_i[11]~input_o ),
	.freq_mod_i_10(\freq_mod_i[10]~input_o ),
	.phi_inc_i_10(\phi_inc_i[10]~input_o ),
	.freq_mod_i_9(\freq_mod_i[9]~input_o ),
	.phi_inc_i_9(\phi_inc_i[9]~input_o ),
	.freq_mod_i_8(\freq_mod_i[8]~input_o ),
	.phi_inc_i_8(\phi_inc_i[8]~input_o ),
	.freq_mod_i_7(\freq_mod_i[7]~input_o ),
	.phi_inc_i_7(\phi_inc_i[7]~input_o ),
	.freq_mod_i_6(\freq_mod_i[6]~input_o ),
	.phi_inc_i_6(\phi_inc_i[6]~input_o ),
	.freq_mod_i_5(\freq_mod_i[5]~input_o ),
	.phi_inc_i_5(\phi_inc_i[5]~input_o ),
	.freq_mod_i_4(\freq_mod_i[4]~input_o ),
	.phi_inc_i_4(\phi_inc_i[4]~input_o ),
	.freq_mod_i_3(\freq_mod_i[3]~input_o ),
	.phi_inc_i_3(\phi_inc_i[3]~input_o ),
	.freq_mod_i_2(\freq_mod_i[2]~input_o ),
	.phi_inc_i_2(\phi_inc_i[2]~input_o ),
	.freq_mod_i_1(\freq_mod_i[1]~input_o ),
	.phi_inc_i_1(\phi_inc_i[1]~input_o ),
	.freq_mod_i_0(\freq_mod_i[0]~input_o ),
	.phi_inc_i_0(\phi_inc_i[0]~input_o ));

assign \clk~input_o  = clk;

assign \reset_n~input_o  = reset_n;

assign \clken~input_o  = clken;

assign \phase_mod_i[0]~input_o  = phase_mod_i[0];

assign \phase_mod_i[1]~input_o  = phase_mod_i[1];

assign \phase_mod_i[2]~input_o  = phase_mod_i[2];

assign \phase_mod_i[3]~input_o  = phase_mod_i[3];

assign \phase_mod_i[4]~input_o  = phase_mod_i[4];

assign \phase_mod_i[5]~input_o  = phase_mod_i[5];

assign \phase_mod_i[6]~input_o  = phase_mod_i[6];

assign \phase_mod_i[7]~input_o  = phase_mod_i[7];

assign \phase_mod_i[8]~input_o  = phase_mod_i[8];

assign \phase_mod_i[9]~input_o  = phase_mod_i[9];

assign \phase_mod_i[10]~input_o  = phase_mod_i[10];

assign \phase_mod_i[11]~input_o  = phase_mod_i[11];

assign \phase_mod_i[12]~input_o  = phase_mod_i[12];

assign \phase_mod_i[15]~input_o  = phase_mod_i[15];

assign \phase_mod_i[13]~input_o  = phase_mod_i[13];

assign \phase_mod_i[14]~input_o  = phase_mod_i[14];

assign \freq_mod_i[16]~input_o  = freq_mod_i[16];

assign \phi_inc_i[16]~input_o  = phi_inc_i[16];

assign \freq_mod_i[17]~input_o  = freq_mod_i[17];

assign \phi_inc_i[17]~input_o  = phi_inc_i[17];

assign \freq_mod_i[18]~input_o  = freq_mod_i[18];

assign \phi_inc_i[18]~input_o  = phi_inc_i[18];

assign \freq_mod_i[19]~input_o  = freq_mod_i[19];

assign \phi_inc_i[19]~input_o  = phi_inc_i[19];

assign \freq_mod_i[20]~input_o  = freq_mod_i[20];

assign \phi_inc_i[20]~input_o  = phi_inc_i[20];

assign \freq_mod_i[21]~input_o  = freq_mod_i[21];

assign \phi_inc_i[21]~input_o  = phi_inc_i[21];

assign \freq_mod_i[22]~input_o  = freq_mod_i[22];

assign \phi_inc_i[22]~input_o  = phi_inc_i[22];

assign \freq_mod_i[23]~input_o  = freq_mod_i[23];

assign \phi_inc_i[23]~input_o  = phi_inc_i[23];

assign \freq_mod_i[24]~input_o  = freq_mod_i[24];

assign \phi_inc_i[24]~input_o  = phi_inc_i[24];

assign \freq_mod_i[25]~input_o  = freq_mod_i[25];

assign \phi_inc_i[25]~input_o  = phi_inc_i[25];

assign \freq_mod_i[26]~input_o  = freq_mod_i[26];

assign \phi_inc_i[26]~input_o  = phi_inc_i[26];

assign \freq_mod_i[27]~input_o  = freq_mod_i[27];

assign \phi_inc_i[27]~input_o  = phi_inc_i[27];

assign \freq_mod_i[28]~input_o  = freq_mod_i[28];

assign \phi_inc_i[28]~input_o  = phi_inc_i[28];

assign \freq_mod_i[31]~input_o  = freq_mod_i[31];

assign \phi_inc_i[31]~input_o  = phi_inc_i[31];

assign \freq_mod_i[15]~input_o  = freq_mod_i[15];

assign \phi_inc_i[15]~input_o  = phi_inc_i[15];

assign \freq_mod_i[29]~input_o  = freq_mod_i[29];

assign \phi_inc_i[29]~input_o  = phi_inc_i[29];

assign \freq_mod_i[30]~input_o  = freq_mod_i[30];

assign \phi_inc_i[30]~input_o  = phi_inc_i[30];

assign \freq_mod_i[14]~input_o  = freq_mod_i[14];

assign \phi_inc_i[14]~input_o  = phi_inc_i[14];

assign \freq_mod_i[13]~input_o  = freq_mod_i[13];

assign \phi_inc_i[13]~input_o  = phi_inc_i[13];

assign \freq_mod_i[12]~input_o  = freq_mod_i[12];

assign \phi_inc_i[12]~input_o  = phi_inc_i[12];

assign \freq_mod_i[11]~input_o  = freq_mod_i[11];

assign \phi_inc_i[11]~input_o  = phi_inc_i[11];

assign \freq_mod_i[10]~input_o  = freq_mod_i[10];

assign \phi_inc_i[10]~input_o  = phi_inc_i[10];

assign \freq_mod_i[9]~input_o  = freq_mod_i[9];

assign \phi_inc_i[9]~input_o  = phi_inc_i[9];

assign \freq_mod_i[8]~input_o  = freq_mod_i[8];

assign \phi_inc_i[8]~input_o  = phi_inc_i[8];

assign \freq_mod_i[7]~input_o  = freq_mod_i[7];

assign \phi_inc_i[7]~input_o  = phi_inc_i[7];

assign \freq_mod_i[6]~input_o  = freq_mod_i[6];

assign \phi_inc_i[6]~input_o  = phi_inc_i[6];

assign \freq_mod_i[5]~input_o  = freq_mod_i[5];

assign \phi_inc_i[5]~input_o  = phi_inc_i[5];

assign \freq_mod_i[4]~input_o  = freq_mod_i[4];

assign \phi_inc_i[4]~input_o  = phi_inc_i[4];

assign \freq_mod_i[3]~input_o  = freq_mod_i[3];

assign \phi_inc_i[3]~input_o  = phi_inc_i[3];

assign \freq_mod_i[2]~input_o  = freq_mod_i[2];

assign \phi_inc_i[2]~input_o  = phi_inc_i[2];

assign \freq_mod_i[1]~input_o  = freq_mod_i[1];

assign \phi_inc_i[1]~input_o  = phi_inc_i[1];

assign \freq_mod_i[0]~input_o  = freq_mod_i[0];

assign \phi_inc_i[0]~input_o  = phi_inc_i[0];

assign fsin_o[0] = \nco_ii_0|ux122|data_out[0]~q ;

assign fsin_o[1] = \nco_ii_0|ux122|data_out[1]~q ;

assign fsin_o[2] = \nco_ii_0|ux122|data_out[2]~q ;

assign fsin_o[3] = \nco_ii_0|ux122|data_out[3]~q ;

assign fsin_o[4] = \nco_ii_0|ux122|data_out[4]~q ;

assign fsin_o[5] = \nco_ii_0|ux122|data_out[5]~q ;

assign fsin_o[6] = \nco_ii_0|ux122|data_out[6]~q ;

assign fsin_o[7] = \nco_ii_0|ux122|data_out[7]~q ;

assign fsin_o[8] = \nco_ii_0|ux122|data_out[8]~q ;

assign fsin_o[9] = \nco_ii_0|ux122|data_out[9]~q ;

assign fsin_o[10] = \nco_ii_0|ux122|data_out[10]~q ;

assign fsin_o[11] = \nco_ii_0|ux122|data_out[11]~q ;

assign fsin_o[12] = \nco_ii_0|ux122|data_out[12]~q ;

assign fsin_o[13] = \nco_ii_0|ux122|data_out[13]~q ;

assign fsin_o[14] = \nco_ii_0|ux122|data_out[14]~q ;

assign fsin_o[15] = \nco_ii_0|ux122|data_out[15]~q ;

assign fsin_o[16] = \nco_ii_0|ux122|data_out[16]~q ;

assign fsin_o[17] = \nco_ii_0|ux122|data_out[17]~q ;

assign fsin_o[18] = \nco_ii_0|ux122|data_out[18]~q ;

assign fsin_o[19] = \nco_ii_0|ux122|data_out[19]~q ;

assign fsin_o[20] = \nco_ii_0|ux122|data_out[20]~q ;

assign fsin_o[21] = \nco_ii_0|ux122|data_out[21]~q ;

assign fsin_o[22] = \nco_ii_0|ux122|data_out[22]~q ;

assign fsin_o[23] = \nco_ii_0|ux122|data_out[23]~q ;

assign out_valid = \nco_ii_0|ux710isdr|data_ready~q ;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cyclonev_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 64'h6666666666666666;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 64'h9696969696969696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cyclonev_lcell_comb \~QIC_CREATED_GND~I (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~QIC_CREATED_GND~I_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~QIC_CREATED_GND~I .extended_lut = "off";
defparam \~QIC_CREATED_GND~I .lut_mask = 64'h0000000000000000;
defparam \~QIC_CREATED_GND~I .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\~QIC_CREATED_GND~I_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3 .lut_mask = 64'hF9F6FFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 .lut_mask = 64'hFF96FFFFFF96FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .lut_mask = 64'h7FFFDFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .lut_mask = 64'h6666666666666666;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .lut_mask = 64'h6666666666666666;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .lut_mask = 64'hDEDEDEDEDEDEDEDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .lut_mask = 64'hEDDEEDDEEDDEEDDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .lut_mask = 64'hDEEDEDDEDEEDEDDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .lut_mask = 64'hEDDEDEEDDEEDEDDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .lut_mask = 64'hBEBEBEBEBEBEBEBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .lut_mask = 64'hBEEBEBBEBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .lut_mask = 64'hBEEBEBBEBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|SQHZ7915_1 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_1 .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|SQHZ7915_2 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_2 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 64'hFDF7FFFFF7FDFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 64'hDFD5FFFFDFD5FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|AMGP4450~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|AMGP4450 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|AMGP4450 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|AMGP4450 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|NJQG9082~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|NJQG9082 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 64'hCF5FFFFFCF5FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .lut_mask = 64'hAFFAAFFAAFFAAFFA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .lut_mask = 64'hBEEBBEEBEBBEEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .lut_mask = 64'hFFFFFFBFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 64'hFFFFFFF6FFFFFFF6;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 64'hD1FFD1FFD1FFD1FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .lut_mask = 64'hF7D5F7D5F7D5F7D5;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .lut_mask = 64'hD8FFFFFFD8FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 64'hEFFFFEFFEFFFFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~5_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 .lut_mask = 64'hFFEFFFFFFFEFFFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 .lut_mask = 64'hBFEFFFFFBFEFFFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 .lut_mask = 64'hFBFEEBBEFBFEEBBE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|comb~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|comb~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|comb~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \nabboc|pzdyqx_impl_inst|comb~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .lut_mask = 64'h6996F9F66996F9F6;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .lut_mask = 64'hDDF5DFFDDDF5DFFD;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 .lut_mask = 64'h6996F9F66996F9F6;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datae(!\altera_internal_jtag~TDIUTAP ),
	.dataf(!\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 .lut_mask = 64'hB1FFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|sdr (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|sdr .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|sdr .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \nabboc|pzdyqx_impl_inst|sdr .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|dr_scan (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|dr_scan .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|dr_scan .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \nabboc|pzdyqx_impl_inst|dr_scan .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|KNOR6738 (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|tdo~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .lut_mask = 64'hFF55FF55FF55FF55;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .lut_mask = 64'h55FFFF5555FFFF55;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .lut_mask = 64'hDD7777DDDD7777DD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .lut_mask = 64'hD77D7DD77DD7D77D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 64'hFFFF6996FFFF6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .lut_mask = 64'hFFFF6996FFFF6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .lut_mask = 64'hFFFF6996FFFF6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|~GND .extended_lut = "off";
defparam \auto_hub|~GND .lut_mask = 64'h0000000000000000;
defparam \auto_hub|~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .shared_arith = "off";

endmodule

module sine_sine_nco_ii_0 (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	data_out_10,
	data_out_11,
	data_out_12,
	data_out_13,
	data_out_14,
	data_out_15,
	data_out_16,
	data_out_17,
	data_out_18,
	data_out_19,
	data_out_20,
	data_out_21,
	data_out_22,
	data_out_23,
	data_ready,
	NJQG9082,
	clk,
	reset_n,
	clken,
	phase_mod_i_0,
	phase_mod_i_1,
	phase_mod_i_2,
	phase_mod_i_3,
	phase_mod_i_4,
	phase_mod_i_5,
	phase_mod_i_6,
	phase_mod_i_7,
	phase_mod_i_8,
	phase_mod_i_9,
	phase_mod_i_10,
	phase_mod_i_11,
	phase_mod_i_12,
	phase_mod_i_15,
	phase_mod_i_13,
	phase_mod_i_14,
	freq_mod_i_16,
	phi_inc_i_16,
	freq_mod_i_17,
	phi_inc_i_17,
	freq_mod_i_18,
	phi_inc_i_18,
	freq_mod_i_19,
	phi_inc_i_19,
	freq_mod_i_20,
	phi_inc_i_20,
	freq_mod_i_21,
	phi_inc_i_21,
	freq_mod_i_22,
	phi_inc_i_22,
	freq_mod_i_23,
	phi_inc_i_23,
	freq_mod_i_24,
	phi_inc_i_24,
	freq_mod_i_25,
	phi_inc_i_25,
	freq_mod_i_26,
	phi_inc_i_26,
	freq_mod_i_27,
	phi_inc_i_27,
	freq_mod_i_28,
	phi_inc_i_28,
	freq_mod_i_31,
	phi_inc_i_31,
	freq_mod_i_15,
	phi_inc_i_15,
	freq_mod_i_29,
	phi_inc_i_29,
	freq_mod_i_30,
	phi_inc_i_30,
	freq_mod_i_14,
	phi_inc_i_14,
	freq_mod_i_13,
	phi_inc_i_13,
	freq_mod_i_12,
	phi_inc_i_12,
	freq_mod_i_11,
	phi_inc_i_11,
	freq_mod_i_10,
	phi_inc_i_10,
	freq_mod_i_9,
	phi_inc_i_9,
	freq_mod_i_8,
	phi_inc_i_8,
	freq_mod_i_7,
	phi_inc_i_7,
	freq_mod_i_6,
	phi_inc_i_6,
	freq_mod_i_5,
	phi_inc_i_5,
	freq_mod_i_4,
	phi_inc_i_4,
	freq_mod_i_3,
	phi_inc_i_3,
	freq_mod_i_2,
	phi_inc_i_2,
	freq_mod_i_1,
	phi_inc_i_1,
	freq_mod_i_0,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
output 	data_out_8;
output 	data_out_9;
output 	data_out_10;
output 	data_out_11;
output 	data_out_12;
output 	data_out_13;
output 	data_out_14;
output 	data_out_15;
output 	data_out_16;
output 	data_out_17;
output 	data_out_18;
output 	data_out_19;
output 	data_out_20;
output 	data_out_21;
output 	data_out_22;
output 	data_out_23;
output 	data_ready;
input 	NJQG9082;
input 	clk;
input 	reset_n;
input 	clken;
input 	phase_mod_i_0;
input 	phase_mod_i_1;
input 	phase_mod_i_2;
input 	phase_mod_i_3;
input 	phase_mod_i_4;
input 	phase_mod_i_5;
input 	phase_mod_i_6;
input 	phase_mod_i_7;
input 	phase_mod_i_8;
input 	phase_mod_i_9;
input 	phase_mod_i_10;
input 	phase_mod_i_11;
input 	phase_mod_i_12;
input 	phase_mod_i_15;
input 	phase_mod_i_13;
input 	phase_mod_i_14;
input 	freq_mod_i_16;
input 	phi_inc_i_16;
input 	freq_mod_i_17;
input 	phi_inc_i_17;
input 	freq_mod_i_18;
input 	phi_inc_i_18;
input 	freq_mod_i_19;
input 	phi_inc_i_19;
input 	freq_mod_i_20;
input 	phi_inc_i_20;
input 	freq_mod_i_21;
input 	phi_inc_i_21;
input 	freq_mod_i_22;
input 	phi_inc_i_22;
input 	freq_mod_i_23;
input 	phi_inc_i_23;
input 	freq_mod_i_24;
input 	phi_inc_i_24;
input 	freq_mod_i_25;
input 	phi_inc_i_25;
input 	freq_mod_i_26;
input 	phi_inc_i_26;
input 	freq_mod_i_27;
input 	phi_inc_i_27;
input 	freq_mod_i_28;
input 	phi_inc_i_28;
input 	freq_mod_i_31;
input 	phi_inc_i_31;
input 	freq_mod_i_15;
input 	phi_inc_i_15;
input 	freq_mod_i_29;
input 	phi_inc_i_29;
input 	freq_mod_i_30;
input 	phi_inc_i_30;
input 	freq_mod_i_14;
input 	phi_inc_i_14;
input 	freq_mod_i_13;
input 	phi_inc_i_13;
input 	freq_mod_i_12;
input 	phi_inc_i_12;
input 	freq_mod_i_11;
input 	phi_inc_i_11;
input 	freq_mod_i_10;
input 	phi_inc_i_10;
input 	freq_mod_i_9;
input 	phi_inc_i_9;
input 	freq_mod_i_8;
input 	phi_inc_i_8;
input 	freq_mod_i_7;
input 	phi_inc_i_7;
input 	freq_mod_i_6;
input 	phi_inc_i_6;
input 	freq_mod_i_5;
input 	phi_inc_i_5;
input 	freq_mod_i_4;
input 	phi_inc_i_4;
input 	freq_mod_i_3;
input 	phi_inc_i_3;
input 	freq_mod_i_2;
input 	phi_inc_i_2;
input 	freq_mod_i_1;
input 	phi_inc_i_1;
input 	freq_mod_i_0;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ux0120|altsyncram_component0|auto_generated|ram_block1a96~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a120~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a144~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a168~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a48~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a72~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a0~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a24~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a97~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a121~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a145~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a169~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a49~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a73~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a1~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a25~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a98~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a122~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a146~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a170~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a50~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a74~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a2~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a26~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a99~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a123~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a147~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a171~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a51~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a75~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a3~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a27~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a100~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a124~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a148~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a172~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a52~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a76~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a4~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a28~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a101~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a125~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a149~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a173~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a53~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a77~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a5~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a29~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a102~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a126~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a150~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a174~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a54~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a78~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a6~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a30~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a103~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a127~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a151~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a175~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a55~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a79~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a7~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a31~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a104~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a128~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a152~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a176~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a56~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a80~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a8~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a32~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a105~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a129~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a153~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a177~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a57~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a81~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a9~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a33~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a106~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a130~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a154~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a178~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a58~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a82~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a10~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a34~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a107~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a131~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a155~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a179~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a59~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a83~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a11~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a35~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a108~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a132~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a156~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a180~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a60~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a84~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a12~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a36~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a109~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a133~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a157~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a181~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a61~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a85~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a13~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a37~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a110~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a134~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a158~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a182~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a62~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a86~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a14~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a38~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a111~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a135~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a159~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a183~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a63~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a87~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a15~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a39~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a112~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a136~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a160~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a184~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a64~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a88~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a16~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a40~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a113~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a137~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a161~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a185~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a65~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a89~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a17~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a41~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a114~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a138~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a162~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a186~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a66~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a90~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a18~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a42~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a115~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a139~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a163~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a187~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a67~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a91~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a19~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a43~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a116~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a140~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a164~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a188~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a68~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a92~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a20~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a44~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a117~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a141~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a165~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a189~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a69~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a93~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a21~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a45~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a118~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a142~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a166~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a190~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a70~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a94~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a22~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a46~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a119~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a143~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a167~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a191~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a71~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a95~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a23~portadataout ;
wire \ux0120|altsyncram_component0|auto_generated|ram_block1a47~portadataout ;
wire \ux009|rom_add[0]~q ;
wire \ux009|rom_add[1]~q ;
wire \ux009|rom_add[2]~q ;
wire \ux009|rom_add[3]~q ;
wire \ux009|rom_add[4]~q ;
wire \ux009|rom_add[5]~q ;
wire \ux009|rom_add[6]~q ;
wire \ux009|rom_add[7]~q ;
wire \ux009|rom_add[8]~q ;
wire \ux009|rom_add[9]~q ;
wire \ux009|rom_add[10]~q ;
wire \ux009|rom_add[11]~q ;
wire \ux009|rom_add[12]~q ;
wire \ux009|rom_add[15]~q ;
wire \ux009|rom_add[13]~q ;
wire \ux009|rom_add[14]~q ;
wire \ux002|dxxpdo[5]~q ;
wire \ux002|dxxpdo[6]~q ;
wire \ux002|dxxpdo[7]~q ;
wire \ux002|dxxpdo[8]~q ;
wire \ux002|dxxpdo[9]~q ;
wire \ux002|dxxpdo[10]~q ;
wire \ux002|dxxpdo[11]~q ;
wire \ux002|dxxpdo[12]~q ;
wire \ux002|dxxpdo[13]~q ;
wire \ux002|dxxpdo[14]~q ;
wire \ux002|dxxpdo[15]~q ;
wire \ux002|dxxpdo[16]~q ;
wire \ux002|dxxpdo[17]~q ;
wire \ux002|dxxpdo[20]~q ;
wire \ux002|dxxpdo[18]~q ;
wire \ux002|dxxpdo[19]~q ;
wire \ux001|dxxrv[3]~q ;
wire \ux001|dxxrv[2]~q ;
wire \ux001|dxxrv[1]~q ;
wire \ux001|dxxrv[0]~q ;
wire \ux0120|altsyncram_component0|auto_generated|out_address_reg_a[2]~q ;
wire \ux0120|altsyncram_component0|auto_generated|out_address_reg_a[0]~q ;
wire \ux0120|altsyncram_component0|auto_generated|out_address_reg_a[1]~q ;
wire \ux122|data_out[12]~3_combout ;
wire \ux004|acc|auto_generated|pipeline_dffe[0]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[1]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[2]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[3]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[4]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[5]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[6]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[7]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[8]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[9]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[10]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[11]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[12]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[15]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[13]~q ;
wire \ux004|acc|auto_generated|pipeline_dffe[14]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[16]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[17]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[18]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[19]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[20]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[21]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[22]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[23]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[24]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[25]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[26]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[27]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[28]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[31]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[15]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[29]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[30]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[14]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[16]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[13]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[17]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[18]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[19]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[20]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[21]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[22]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[23]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[24]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[25]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[26]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[27]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[28]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[31]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[15]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[12]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[29]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[30]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[14]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[11]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[13]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[12]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[11]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[10]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[9]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[8]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[7]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[6]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[5]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[4]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[3]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[2]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[1]~q ;
wire \ux003|acc|auto_generated|pipeline_dffe[0]~q ;


sine_asj_altqmcpipe ux000(
	.data_out_12(\ux122|data_out[12]~3_combout ),
	.pipeline_dffe_16(\ux000|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\ux000|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\ux000|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_19(\ux000|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_20(\ux000|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_21(\ux000|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_22(\ux000|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_23(\ux000|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_24(\ux000|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_25(\ux000|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_26(\ux000|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_27(\ux000|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_28(\ux000|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_31(\ux000|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_15(\ux000|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_29(\ux000|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_30(\ux000|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_14(\ux000|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_161(\ux003|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_13(\ux000|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_171(\ux003|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_181(\ux003|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_191(\ux003|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_201(\ux003|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_211(\ux003|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_221(\ux003|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_231(\ux003|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_241(\ux003|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_251(\ux003|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_261(\ux003|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_271(\ux003|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_281(\ux003|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_311(\ux003|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_151(\ux003|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\ux000|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_291(\ux003|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_301(\ux003|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_141(\ux003|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_11(\ux000|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_131(\ux003|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_121(\ux003|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_111(\ux003|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\ux003|acc|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_9(\ux003|acc|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\ux003|acc|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\ux003|acc|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_6(\ux003|acc|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\ux003|acc|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\ux003|acc|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\ux003|acc|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\ux003|acc|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_1(\ux003|acc|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_0(\ux003|acc|auto_generated|pipeline_dffe[0]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

sine_asj_nco_fxx ux003(
	.pipeline_dffe_16(\ux003|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\ux003|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\ux003|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_19(\ux003|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_20(\ux003|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_21(\ux003|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_22(\ux003|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_23(\ux003|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_24(\ux003|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_25(\ux003|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_26(\ux003|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_27(\ux003|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_28(\ux003|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_31(\ux003|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_15(\ux003|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_29(\ux003|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_30(\ux003|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_14(\ux003|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\ux003|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_12(\ux003|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\ux003|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\ux003|acc|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_9(\ux003|acc|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\ux003|acc|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\ux003|acc|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_6(\ux003|acc|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\ux003|acc|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\ux003|acc|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\ux003|acc|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\ux003|acc|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_1(\ux003|acc|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_0(\ux003|acc|auto_generated|pipeline_dffe[0]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken),
	.freq_mod_i_16(freq_mod_i_16),
	.phi_inc_i_16(phi_inc_i_16),
	.freq_mod_i_17(freq_mod_i_17),
	.phi_inc_i_17(phi_inc_i_17),
	.freq_mod_i_18(freq_mod_i_18),
	.phi_inc_i_18(phi_inc_i_18),
	.freq_mod_i_19(freq_mod_i_19),
	.phi_inc_i_19(phi_inc_i_19),
	.freq_mod_i_20(freq_mod_i_20),
	.phi_inc_i_20(phi_inc_i_20),
	.freq_mod_i_21(freq_mod_i_21),
	.phi_inc_i_21(phi_inc_i_21),
	.freq_mod_i_22(freq_mod_i_22),
	.phi_inc_i_22(phi_inc_i_22),
	.freq_mod_i_23(freq_mod_i_23),
	.phi_inc_i_23(phi_inc_i_23),
	.freq_mod_i_24(freq_mod_i_24),
	.phi_inc_i_24(phi_inc_i_24),
	.freq_mod_i_25(freq_mod_i_25),
	.phi_inc_i_25(phi_inc_i_25),
	.freq_mod_i_26(freq_mod_i_26),
	.phi_inc_i_26(phi_inc_i_26),
	.freq_mod_i_27(freq_mod_i_27),
	.phi_inc_i_27(phi_inc_i_27),
	.freq_mod_i_28(freq_mod_i_28),
	.phi_inc_i_28(phi_inc_i_28),
	.freq_mod_i_31(freq_mod_i_31),
	.phi_inc_i_31(phi_inc_i_31),
	.freq_mod_i_15(freq_mod_i_15),
	.phi_inc_i_15(phi_inc_i_15),
	.freq_mod_i_29(freq_mod_i_29),
	.phi_inc_i_29(phi_inc_i_29),
	.freq_mod_i_30(freq_mod_i_30),
	.phi_inc_i_30(phi_inc_i_30),
	.freq_mod_i_14(freq_mod_i_14),
	.phi_inc_i_14(phi_inc_i_14),
	.freq_mod_i_13(freq_mod_i_13),
	.phi_inc_i_13(phi_inc_i_13),
	.freq_mod_i_12(freq_mod_i_12),
	.phi_inc_i_12(phi_inc_i_12),
	.freq_mod_i_11(freq_mod_i_11),
	.phi_inc_i_11(phi_inc_i_11),
	.freq_mod_i_10(freq_mod_i_10),
	.phi_inc_i_10(phi_inc_i_10),
	.freq_mod_i_9(freq_mod_i_9),
	.phi_inc_i_9(phi_inc_i_9),
	.freq_mod_i_8(freq_mod_i_8),
	.phi_inc_i_8(phi_inc_i_8),
	.freq_mod_i_7(freq_mod_i_7),
	.phi_inc_i_7(phi_inc_i_7),
	.freq_mod_i_6(freq_mod_i_6),
	.phi_inc_i_6(phi_inc_i_6),
	.freq_mod_i_5(freq_mod_i_5),
	.phi_inc_i_5(phi_inc_i_5),
	.freq_mod_i_4(freq_mod_i_4),
	.phi_inc_i_4(phi_inc_i_4),
	.freq_mod_i_3(freq_mod_i_3),
	.phi_inc_i_3(phi_inc_i_3),
	.freq_mod_i_2(freq_mod_i_2),
	.phi_inc_i_2(phi_inc_i_2),
	.freq_mod_i_1(freq_mod_i_1),
	.phi_inc_i_1(phi_inc_i_1),
	.freq_mod_i_0(freq_mod_i_0),
	.phi_inc_i_0(phi_inc_i_0));

sine_asj_nco_pxx ux004(
	.dxxpdo_5(\ux002|dxxpdo[5]~q ),
	.dxxpdo_6(\ux002|dxxpdo[6]~q ),
	.dxxpdo_7(\ux002|dxxpdo[7]~q ),
	.dxxpdo_8(\ux002|dxxpdo[8]~q ),
	.dxxpdo_9(\ux002|dxxpdo[9]~q ),
	.dxxpdo_10(\ux002|dxxpdo[10]~q ),
	.dxxpdo_11(\ux002|dxxpdo[11]~q ),
	.dxxpdo_12(\ux002|dxxpdo[12]~q ),
	.dxxpdo_13(\ux002|dxxpdo[13]~q ),
	.dxxpdo_14(\ux002|dxxpdo[14]~q ),
	.dxxpdo_15(\ux002|dxxpdo[15]~q ),
	.dxxpdo_16(\ux002|dxxpdo[16]~q ),
	.dxxpdo_17(\ux002|dxxpdo[17]~q ),
	.dxxpdo_20(\ux002|dxxpdo[20]~q ),
	.dxxpdo_18(\ux002|dxxpdo[18]~q ),
	.dxxpdo_19(\ux002|dxxpdo[19]~q ),
	.data_out_12(\ux122|data_out[12]~3_combout ),
	.pipeline_dffe_0(\ux004|acc|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\ux004|acc|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\ux004|acc|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\ux004|acc|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\ux004|acc|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\ux004|acc|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\ux004|acc|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\ux004|acc|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\ux004|acc|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\ux004|acc|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\ux004|acc|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\ux004|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\ux004|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_15(\ux004|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_13(\ux004|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\ux004|acc|auto_generated|pipeline_dffe[14]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken),
	.phase_mod_i_0(phase_mod_i_0),
	.phase_mod_i_1(phase_mod_i_1),
	.phase_mod_i_2(phase_mod_i_2),
	.phase_mod_i_3(phase_mod_i_3),
	.phase_mod_i_4(phase_mod_i_4),
	.phase_mod_i_5(phase_mod_i_5),
	.phase_mod_i_6(phase_mod_i_6),
	.phase_mod_i_7(phase_mod_i_7),
	.phase_mod_i_8(phase_mod_i_8),
	.phase_mod_i_9(phase_mod_i_9),
	.phase_mod_i_10(phase_mod_i_10),
	.phase_mod_i_11(phase_mod_i_11),
	.phase_mod_i_12(phase_mod_i_12),
	.phase_mod_i_15(phase_mod_i_15),
	.phase_mod_i_13(phase_mod_i_13),
	.phase_mod_i_14(phase_mod_i_14));

sine_asj_dxx ux002(
	.dxxpdo_5(\ux002|dxxpdo[5]~q ),
	.dxxpdo_6(\ux002|dxxpdo[6]~q ),
	.dxxpdo_7(\ux002|dxxpdo[7]~q ),
	.dxxpdo_8(\ux002|dxxpdo[8]~q ),
	.dxxpdo_9(\ux002|dxxpdo[9]~q ),
	.dxxpdo_10(\ux002|dxxpdo[10]~q ),
	.dxxpdo_11(\ux002|dxxpdo[11]~q ),
	.dxxpdo_12(\ux002|dxxpdo[12]~q ),
	.dxxpdo_13(\ux002|dxxpdo[13]~q ),
	.dxxpdo_14(\ux002|dxxpdo[14]~q ),
	.dxxpdo_15(\ux002|dxxpdo[15]~q ),
	.dxxpdo_16(\ux002|dxxpdo[16]~q ),
	.dxxpdo_17(\ux002|dxxpdo[17]~q ),
	.dxxpdo_20(\ux002|dxxpdo[20]~q ),
	.dxxpdo_18(\ux002|dxxpdo[18]~q ),
	.dxxpdo_19(\ux002|dxxpdo[19]~q ),
	.dxxrv_3(\ux001|dxxrv[3]~q ),
	.dxxrv_2(\ux001|dxxrv[2]~q ),
	.dxxrv_1(\ux001|dxxrv[1]~q ),
	.dxxrv_0(\ux001|dxxrv[0]~q ),
	.data_out_12(\ux122|data_out[12]~3_combout ),
	.pipeline_dffe_16(\ux000|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\ux000|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_18(\ux000|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_19(\ux000|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_20(\ux000|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_21(\ux000|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_22(\ux000|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_23(\ux000|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_24(\ux000|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_25(\ux000|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_26(\ux000|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_27(\ux000|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_28(\ux000|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_31(\ux000|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_15(\ux000|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_29(\ux000|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_30(\ux000|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_14(\ux000|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\ux000|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_12(\ux000|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\ux000|acc|auto_generated|pipeline_dffe[11]~q ),
	.NJQG9082(NJQG9082),
	.clk(clk),
	.reset_n(reset_n));

sine_asj_dxx_g ux001(
	.dxxrv_3(\ux001|dxxrv[3]~q ),
	.dxxrv_2(\ux001|dxxrv[2]~q ),
	.dxxrv_1(\ux001|dxxrv[1]~q ),
	.dxxrv_0(\ux001|dxxrv[0]~q ),
	.data_out_12(\ux122|data_out[12]~3_combout ),
	.clk(clk),
	.reset_n(reset_n));

sine_asj_nco_as_m_cen ux0120(
	.ram_block1a96(\ux0120|altsyncram_component0|auto_generated|ram_block1a96~portadataout ),
	.ram_block1a120(\ux0120|altsyncram_component0|auto_generated|ram_block1a120~portadataout ),
	.ram_block1a144(\ux0120|altsyncram_component0|auto_generated|ram_block1a144~portadataout ),
	.ram_block1a168(\ux0120|altsyncram_component0|auto_generated|ram_block1a168~portadataout ),
	.ram_block1a48(\ux0120|altsyncram_component0|auto_generated|ram_block1a48~portadataout ),
	.ram_block1a72(\ux0120|altsyncram_component0|auto_generated|ram_block1a72~portadataout ),
	.ram_block1a0(\ux0120|altsyncram_component0|auto_generated|ram_block1a0~portadataout ),
	.ram_block1a24(\ux0120|altsyncram_component0|auto_generated|ram_block1a24~portadataout ),
	.ram_block1a97(\ux0120|altsyncram_component0|auto_generated|ram_block1a97~portadataout ),
	.ram_block1a121(\ux0120|altsyncram_component0|auto_generated|ram_block1a121~portadataout ),
	.ram_block1a145(\ux0120|altsyncram_component0|auto_generated|ram_block1a145~portadataout ),
	.ram_block1a169(\ux0120|altsyncram_component0|auto_generated|ram_block1a169~portadataout ),
	.ram_block1a49(\ux0120|altsyncram_component0|auto_generated|ram_block1a49~portadataout ),
	.ram_block1a73(\ux0120|altsyncram_component0|auto_generated|ram_block1a73~portadataout ),
	.ram_block1a1(\ux0120|altsyncram_component0|auto_generated|ram_block1a1~portadataout ),
	.ram_block1a25(\ux0120|altsyncram_component0|auto_generated|ram_block1a25~portadataout ),
	.ram_block1a98(\ux0120|altsyncram_component0|auto_generated|ram_block1a98~portadataout ),
	.ram_block1a122(\ux0120|altsyncram_component0|auto_generated|ram_block1a122~portadataout ),
	.ram_block1a146(\ux0120|altsyncram_component0|auto_generated|ram_block1a146~portadataout ),
	.ram_block1a170(\ux0120|altsyncram_component0|auto_generated|ram_block1a170~portadataout ),
	.ram_block1a50(\ux0120|altsyncram_component0|auto_generated|ram_block1a50~portadataout ),
	.ram_block1a74(\ux0120|altsyncram_component0|auto_generated|ram_block1a74~portadataout ),
	.ram_block1a2(\ux0120|altsyncram_component0|auto_generated|ram_block1a2~portadataout ),
	.ram_block1a26(\ux0120|altsyncram_component0|auto_generated|ram_block1a26~portadataout ),
	.ram_block1a99(\ux0120|altsyncram_component0|auto_generated|ram_block1a99~portadataout ),
	.ram_block1a123(\ux0120|altsyncram_component0|auto_generated|ram_block1a123~portadataout ),
	.ram_block1a147(\ux0120|altsyncram_component0|auto_generated|ram_block1a147~portadataout ),
	.ram_block1a171(\ux0120|altsyncram_component0|auto_generated|ram_block1a171~portadataout ),
	.ram_block1a51(\ux0120|altsyncram_component0|auto_generated|ram_block1a51~portadataout ),
	.ram_block1a75(\ux0120|altsyncram_component0|auto_generated|ram_block1a75~portadataout ),
	.ram_block1a3(\ux0120|altsyncram_component0|auto_generated|ram_block1a3~portadataout ),
	.ram_block1a27(\ux0120|altsyncram_component0|auto_generated|ram_block1a27~portadataout ),
	.ram_block1a100(\ux0120|altsyncram_component0|auto_generated|ram_block1a100~portadataout ),
	.ram_block1a124(\ux0120|altsyncram_component0|auto_generated|ram_block1a124~portadataout ),
	.ram_block1a148(\ux0120|altsyncram_component0|auto_generated|ram_block1a148~portadataout ),
	.ram_block1a172(\ux0120|altsyncram_component0|auto_generated|ram_block1a172~portadataout ),
	.ram_block1a52(\ux0120|altsyncram_component0|auto_generated|ram_block1a52~portadataout ),
	.ram_block1a76(\ux0120|altsyncram_component0|auto_generated|ram_block1a76~portadataout ),
	.ram_block1a4(\ux0120|altsyncram_component0|auto_generated|ram_block1a4~portadataout ),
	.ram_block1a28(\ux0120|altsyncram_component0|auto_generated|ram_block1a28~portadataout ),
	.ram_block1a101(\ux0120|altsyncram_component0|auto_generated|ram_block1a101~portadataout ),
	.ram_block1a125(\ux0120|altsyncram_component0|auto_generated|ram_block1a125~portadataout ),
	.ram_block1a149(\ux0120|altsyncram_component0|auto_generated|ram_block1a149~portadataout ),
	.ram_block1a173(\ux0120|altsyncram_component0|auto_generated|ram_block1a173~portadataout ),
	.ram_block1a53(\ux0120|altsyncram_component0|auto_generated|ram_block1a53~portadataout ),
	.ram_block1a77(\ux0120|altsyncram_component0|auto_generated|ram_block1a77~portadataout ),
	.ram_block1a5(\ux0120|altsyncram_component0|auto_generated|ram_block1a5~portadataout ),
	.ram_block1a29(\ux0120|altsyncram_component0|auto_generated|ram_block1a29~portadataout ),
	.ram_block1a102(\ux0120|altsyncram_component0|auto_generated|ram_block1a102~portadataout ),
	.ram_block1a126(\ux0120|altsyncram_component0|auto_generated|ram_block1a126~portadataout ),
	.ram_block1a150(\ux0120|altsyncram_component0|auto_generated|ram_block1a150~portadataout ),
	.ram_block1a174(\ux0120|altsyncram_component0|auto_generated|ram_block1a174~portadataout ),
	.ram_block1a54(\ux0120|altsyncram_component0|auto_generated|ram_block1a54~portadataout ),
	.ram_block1a78(\ux0120|altsyncram_component0|auto_generated|ram_block1a78~portadataout ),
	.ram_block1a6(\ux0120|altsyncram_component0|auto_generated|ram_block1a6~portadataout ),
	.ram_block1a30(\ux0120|altsyncram_component0|auto_generated|ram_block1a30~portadataout ),
	.ram_block1a103(\ux0120|altsyncram_component0|auto_generated|ram_block1a103~portadataout ),
	.ram_block1a127(\ux0120|altsyncram_component0|auto_generated|ram_block1a127~portadataout ),
	.ram_block1a151(\ux0120|altsyncram_component0|auto_generated|ram_block1a151~portadataout ),
	.ram_block1a175(\ux0120|altsyncram_component0|auto_generated|ram_block1a175~portadataout ),
	.ram_block1a55(\ux0120|altsyncram_component0|auto_generated|ram_block1a55~portadataout ),
	.ram_block1a79(\ux0120|altsyncram_component0|auto_generated|ram_block1a79~portadataout ),
	.ram_block1a7(\ux0120|altsyncram_component0|auto_generated|ram_block1a7~portadataout ),
	.ram_block1a31(\ux0120|altsyncram_component0|auto_generated|ram_block1a31~portadataout ),
	.ram_block1a104(\ux0120|altsyncram_component0|auto_generated|ram_block1a104~portadataout ),
	.ram_block1a128(\ux0120|altsyncram_component0|auto_generated|ram_block1a128~portadataout ),
	.ram_block1a152(\ux0120|altsyncram_component0|auto_generated|ram_block1a152~portadataout ),
	.ram_block1a176(\ux0120|altsyncram_component0|auto_generated|ram_block1a176~portadataout ),
	.ram_block1a56(\ux0120|altsyncram_component0|auto_generated|ram_block1a56~portadataout ),
	.ram_block1a80(\ux0120|altsyncram_component0|auto_generated|ram_block1a80~portadataout ),
	.ram_block1a8(\ux0120|altsyncram_component0|auto_generated|ram_block1a8~portadataout ),
	.ram_block1a32(\ux0120|altsyncram_component0|auto_generated|ram_block1a32~portadataout ),
	.ram_block1a105(\ux0120|altsyncram_component0|auto_generated|ram_block1a105~portadataout ),
	.ram_block1a129(\ux0120|altsyncram_component0|auto_generated|ram_block1a129~portadataout ),
	.ram_block1a153(\ux0120|altsyncram_component0|auto_generated|ram_block1a153~portadataout ),
	.ram_block1a177(\ux0120|altsyncram_component0|auto_generated|ram_block1a177~portadataout ),
	.ram_block1a57(\ux0120|altsyncram_component0|auto_generated|ram_block1a57~portadataout ),
	.ram_block1a81(\ux0120|altsyncram_component0|auto_generated|ram_block1a81~portadataout ),
	.ram_block1a9(\ux0120|altsyncram_component0|auto_generated|ram_block1a9~portadataout ),
	.ram_block1a33(\ux0120|altsyncram_component0|auto_generated|ram_block1a33~portadataout ),
	.ram_block1a106(\ux0120|altsyncram_component0|auto_generated|ram_block1a106~portadataout ),
	.ram_block1a130(\ux0120|altsyncram_component0|auto_generated|ram_block1a130~portadataout ),
	.ram_block1a154(\ux0120|altsyncram_component0|auto_generated|ram_block1a154~portadataout ),
	.ram_block1a178(\ux0120|altsyncram_component0|auto_generated|ram_block1a178~portadataout ),
	.ram_block1a58(\ux0120|altsyncram_component0|auto_generated|ram_block1a58~portadataout ),
	.ram_block1a82(\ux0120|altsyncram_component0|auto_generated|ram_block1a82~portadataout ),
	.ram_block1a10(\ux0120|altsyncram_component0|auto_generated|ram_block1a10~portadataout ),
	.ram_block1a34(\ux0120|altsyncram_component0|auto_generated|ram_block1a34~portadataout ),
	.ram_block1a107(\ux0120|altsyncram_component0|auto_generated|ram_block1a107~portadataout ),
	.ram_block1a131(\ux0120|altsyncram_component0|auto_generated|ram_block1a131~portadataout ),
	.ram_block1a155(\ux0120|altsyncram_component0|auto_generated|ram_block1a155~portadataout ),
	.ram_block1a179(\ux0120|altsyncram_component0|auto_generated|ram_block1a179~portadataout ),
	.ram_block1a59(\ux0120|altsyncram_component0|auto_generated|ram_block1a59~portadataout ),
	.ram_block1a83(\ux0120|altsyncram_component0|auto_generated|ram_block1a83~portadataout ),
	.ram_block1a11(\ux0120|altsyncram_component0|auto_generated|ram_block1a11~portadataout ),
	.ram_block1a35(\ux0120|altsyncram_component0|auto_generated|ram_block1a35~portadataout ),
	.ram_block1a108(\ux0120|altsyncram_component0|auto_generated|ram_block1a108~portadataout ),
	.ram_block1a132(\ux0120|altsyncram_component0|auto_generated|ram_block1a132~portadataout ),
	.ram_block1a156(\ux0120|altsyncram_component0|auto_generated|ram_block1a156~portadataout ),
	.ram_block1a180(\ux0120|altsyncram_component0|auto_generated|ram_block1a180~portadataout ),
	.ram_block1a60(\ux0120|altsyncram_component0|auto_generated|ram_block1a60~portadataout ),
	.ram_block1a84(\ux0120|altsyncram_component0|auto_generated|ram_block1a84~portadataout ),
	.ram_block1a12(\ux0120|altsyncram_component0|auto_generated|ram_block1a12~portadataout ),
	.ram_block1a36(\ux0120|altsyncram_component0|auto_generated|ram_block1a36~portadataout ),
	.ram_block1a109(\ux0120|altsyncram_component0|auto_generated|ram_block1a109~portadataout ),
	.ram_block1a133(\ux0120|altsyncram_component0|auto_generated|ram_block1a133~portadataout ),
	.ram_block1a157(\ux0120|altsyncram_component0|auto_generated|ram_block1a157~portadataout ),
	.ram_block1a181(\ux0120|altsyncram_component0|auto_generated|ram_block1a181~portadataout ),
	.ram_block1a61(\ux0120|altsyncram_component0|auto_generated|ram_block1a61~portadataout ),
	.ram_block1a85(\ux0120|altsyncram_component0|auto_generated|ram_block1a85~portadataout ),
	.ram_block1a13(\ux0120|altsyncram_component0|auto_generated|ram_block1a13~portadataout ),
	.ram_block1a37(\ux0120|altsyncram_component0|auto_generated|ram_block1a37~portadataout ),
	.ram_block1a110(\ux0120|altsyncram_component0|auto_generated|ram_block1a110~portadataout ),
	.ram_block1a134(\ux0120|altsyncram_component0|auto_generated|ram_block1a134~portadataout ),
	.ram_block1a158(\ux0120|altsyncram_component0|auto_generated|ram_block1a158~portadataout ),
	.ram_block1a182(\ux0120|altsyncram_component0|auto_generated|ram_block1a182~portadataout ),
	.ram_block1a62(\ux0120|altsyncram_component0|auto_generated|ram_block1a62~portadataout ),
	.ram_block1a86(\ux0120|altsyncram_component0|auto_generated|ram_block1a86~portadataout ),
	.ram_block1a14(\ux0120|altsyncram_component0|auto_generated|ram_block1a14~portadataout ),
	.ram_block1a38(\ux0120|altsyncram_component0|auto_generated|ram_block1a38~portadataout ),
	.ram_block1a111(\ux0120|altsyncram_component0|auto_generated|ram_block1a111~portadataout ),
	.ram_block1a135(\ux0120|altsyncram_component0|auto_generated|ram_block1a135~portadataout ),
	.ram_block1a159(\ux0120|altsyncram_component0|auto_generated|ram_block1a159~portadataout ),
	.ram_block1a183(\ux0120|altsyncram_component0|auto_generated|ram_block1a183~portadataout ),
	.ram_block1a63(\ux0120|altsyncram_component0|auto_generated|ram_block1a63~portadataout ),
	.ram_block1a87(\ux0120|altsyncram_component0|auto_generated|ram_block1a87~portadataout ),
	.ram_block1a15(\ux0120|altsyncram_component0|auto_generated|ram_block1a15~portadataout ),
	.ram_block1a39(\ux0120|altsyncram_component0|auto_generated|ram_block1a39~portadataout ),
	.ram_block1a112(\ux0120|altsyncram_component0|auto_generated|ram_block1a112~portadataout ),
	.ram_block1a136(\ux0120|altsyncram_component0|auto_generated|ram_block1a136~portadataout ),
	.ram_block1a160(\ux0120|altsyncram_component0|auto_generated|ram_block1a160~portadataout ),
	.ram_block1a184(\ux0120|altsyncram_component0|auto_generated|ram_block1a184~portadataout ),
	.ram_block1a64(\ux0120|altsyncram_component0|auto_generated|ram_block1a64~portadataout ),
	.ram_block1a88(\ux0120|altsyncram_component0|auto_generated|ram_block1a88~portadataout ),
	.ram_block1a16(\ux0120|altsyncram_component0|auto_generated|ram_block1a16~portadataout ),
	.ram_block1a40(\ux0120|altsyncram_component0|auto_generated|ram_block1a40~portadataout ),
	.ram_block1a113(\ux0120|altsyncram_component0|auto_generated|ram_block1a113~portadataout ),
	.ram_block1a137(\ux0120|altsyncram_component0|auto_generated|ram_block1a137~portadataout ),
	.ram_block1a161(\ux0120|altsyncram_component0|auto_generated|ram_block1a161~portadataout ),
	.ram_block1a185(\ux0120|altsyncram_component0|auto_generated|ram_block1a185~portadataout ),
	.ram_block1a65(\ux0120|altsyncram_component0|auto_generated|ram_block1a65~portadataout ),
	.ram_block1a89(\ux0120|altsyncram_component0|auto_generated|ram_block1a89~portadataout ),
	.ram_block1a17(\ux0120|altsyncram_component0|auto_generated|ram_block1a17~portadataout ),
	.ram_block1a41(\ux0120|altsyncram_component0|auto_generated|ram_block1a41~portadataout ),
	.ram_block1a114(\ux0120|altsyncram_component0|auto_generated|ram_block1a114~portadataout ),
	.ram_block1a138(\ux0120|altsyncram_component0|auto_generated|ram_block1a138~portadataout ),
	.ram_block1a162(\ux0120|altsyncram_component0|auto_generated|ram_block1a162~portadataout ),
	.ram_block1a186(\ux0120|altsyncram_component0|auto_generated|ram_block1a186~portadataout ),
	.ram_block1a66(\ux0120|altsyncram_component0|auto_generated|ram_block1a66~portadataout ),
	.ram_block1a90(\ux0120|altsyncram_component0|auto_generated|ram_block1a90~portadataout ),
	.ram_block1a18(\ux0120|altsyncram_component0|auto_generated|ram_block1a18~portadataout ),
	.ram_block1a42(\ux0120|altsyncram_component0|auto_generated|ram_block1a42~portadataout ),
	.ram_block1a115(\ux0120|altsyncram_component0|auto_generated|ram_block1a115~portadataout ),
	.ram_block1a139(\ux0120|altsyncram_component0|auto_generated|ram_block1a139~portadataout ),
	.ram_block1a163(\ux0120|altsyncram_component0|auto_generated|ram_block1a163~portadataout ),
	.ram_block1a187(\ux0120|altsyncram_component0|auto_generated|ram_block1a187~portadataout ),
	.ram_block1a67(\ux0120|altsyncram_component0|auto_generated|ram_block1a67~portadataout ),
	.ram_block1a91(\ux0120|altsyncram_component0|auto_generated|ram_block1a91~portadataout ),
	.ram_block1a19(\ux0120|altsyncram_component0|auto_generated|ram_block1a19~portadataout ),
	.ram_block1a43(\ux0120|altsyncram_component0|auto_generated|ram_block1a43~portadataout ),
	.ram_block1a116(\ux0120|altsyncram_component0|auto_generated|ram_block1a116~portadataout ),
	.ram_block1a140(\ux0120|altsyncram_component0|auto_generated|ram_block1a140~portadataout ),
	.ram_block1a164(\ux0120|altsyncram_component0|auto_generated|ram_block1a164~portadataout ),
	.ram_block1a188(\ux0120|altsyncram_component0|auto_generated|ram_block1a188~portadataout ),
	.ram_block1a68(\ux0120|altsyncram_component0|auto_generated|ram_block1a68~portadataout ),
	.ram_block1a92(\ux0120|altsyncram_component0|auto_generated|ram_block1a92~portadataout ),
	.ram_block1a20(\ux0120|altsyncram_component0|auto_generated|ram_block1a20~portadataout ),
	.ram_block1a44(\ux0120|altsyncram_component0|auto_generated|ram_block1a44~portadataout ),
	.ram_block1a117(\ux0120|altsyncram_component0|auto_generated|ram_block1a117~portadataout ),
	.ram_block1a141(\ux0120|altsyncram_component0|auto_generated|ram_block1a141~portadataout ),
	.ram_block1a165(\ux0120|altsyncram_component0|auto_generated|ram_block1a165~portadataout ),
	.ram_block1a189(\ux0120|altsyncram_component0|auto_generated|ram_block1a189~portadataout ),
	.ram_block1a69(\ux0120|altsyncram_component0|auto_generated|ram_block1a69~portadataout ),
	.ram_block1a93(\ux0120|altsyncram_component0|auto_generated|ram_block1a93~portadataout ),
	.ram_block1a21(\ux0120|altsyncram_component0|auto_generated|ram_block1a21~portadataout ),
	.ram_block1a45(\ux0120|altsyncram_component0|auto_generated|ram_block1a45~portadataout ),
	.ram_block1a118(\ux0120|altsyncram_component0|auto_generated|ram_block1a118~portadataout ),
	.ram_block1a142(\ux0120|altsyncram_component0|auto_generated|ram_block1a142~portadataout ),
	.ram_block1a166(\ux0120|altsyncram_component0|auto_generated|ram_block1a166~portadataout ),
	.ram_block1a190(\ux0120|altsyncram_component0|auto_generated|ram_block1a190~portadataout ),
	.ram_block1a70(\ux0120|altsyncram_component0|auto_generated|ram_block1a70~portadataout ),
	.ram_block1a94(\ux0120|altsyncram_component0|auto_generated|ram_block1a94~portadataout ),
	.ram_block1a22(\ux0120|altsyncram_component0|auto_generated|ram_block1a22~portadataout ),
	.ram_block1a46(\ux0120|altsyncram_component0|auto_generated|ram_block1a46~portadataout ),
	.ram_block1a119(\ux0120|altsyncram_component0|auto_generated|ram_block1a119~portadataout ),
	.ram_block1a143(\ux0120|altsyncram_component0|auto_generated|ram_block1a143~portadataout ),
	.ram_block1a167(\ux0120|altsyncram_component0|auto_generated|ram_block1a167~portadataout ),
	.ram_block1a191(\ux0120|altsyncram_component0|auto_generated|ram_block1a191~portadataout ),
	.ram_block1a71(\ux0120|altsyncram_component0|auto_generated|ram_block1a71~portadataout ),
	.ram_block1a95(\ux0120|altsyncram_component0|auto_generated|ram_block1a95~portadataout ),
	.ram_block1a23(\ux0120|altsyncram_component0|auto_generated|ram_block1a23~portadataout ),
	.ram_block1a47(\ux0120|altsyncram_component0|auto_generated|ram_block1a47~portadataout ),
	.rom_add_0(\ux009|rom_add[0]~q ),
	.rom_add_1(\ux009|rom_add[1]~q ),
	.rom_add_2(\ux009|rom_add[2]~q ),
	.rom_add_3(\ux009|rom_add[3]~q ),
	.rom_add_4(\ux009|rom_add[4]~q ),
	.rom_add_5(\ux009|rom_add[5]~q ),
	.rom_add_6(\ux009|rom_add[6]~q ),
	.rom_add_7(\ux009|rom_add[7]~q ),
	.rom_add_8(\ux009|rom_add[8]~q ),
	.rom_add_9(\ux009|rom_add[9]~q ),
	.rom_add_10(\ux009|rom_add[10]~q ),
	.rom_add_11(\ux009|rom_add[11]~q ),
	.rom_add_12(\ux009|rom_add[12]~q ),
	.rom_add_15(\ux009|rom_add[15]~q ),
	.rom_add_13(\ux009|rom_add[13]~q ),
	.rom_add_14(\ux009|rom_add[14]~q ),
	.out_address_reg_a_2(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[2]~q ),
	.out_address_reg_a_0(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[0]~q ),
	.out_address_reg_a_1(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[1]~q ),
	.clk(clk),
	.clken(clken));

sine_asj_gal ux009(
	.rom_add_0(\ux009|rom_add[0]~q ),
	.rom_add_1(\ux009|rom_add[1]~q ),
	.rom_add_2(\ux009|rom_add[2]~q ),
	.rom_add_3(\ux009|rom_add[3]~q ),
	.rom_add_4(\ux009|rom_add[4]~q ),
	.rom_add_5(\ux009|rom_add[5]~q ),
	.rom_add_6(\ux009|rom_add[6]~q ),
	.rom_add_7(\ux009|rom_add[7]~q ),
	.rom_add_8(\ux009|rom_add[8]~q ),
	.rom_add_9(\ux009|rom_add[9]~q ),
	.rom_add_10(\ux009|rom_add[10]~q ),
	.rom_add_11(\ux009|rom_add[11]~q ),
	.rom_add_12(\ux009|rom_add[12]~q ),
	.rom_add_15(\ux009|rom_add[15]~q ),
	.rom_add_13(\ux009|rom_add[13]~q ),
	.rom_add_14(\ux009|rom_add[14]~q ),
	.data_out_12(\ux122|data_out[12]~3_combout ),
	.pipeline_dffe_0(\ux004|acc|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\ux004|acc|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\ux004|acc|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\ux004|acc|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\ux004|acc|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\ux004|acc|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\ux004|acc|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\ux004|acc|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\ux004|acc|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\ux004|acc|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\ux004|acc|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\ux004|acc|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\ux004|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_15(\ux004|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_13(\ux004|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\ux004|acc|auto_generated|pipeline_dffe[14]~q ),
	.clk(clk),
	.reset_n(reset_n));

sine_asj_nco_isdr ux710isdr(
	.data_ready1(data_ready),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

sine_asj_nco_mob_rw ux122(
	.data_out_0(data_out_0),
	.data_out_1(data_out_1),
	.data_out_2(data_out_2),
	.data_out_3(data_out_3),
	.data_out_4(data_out_4),
	.data_out_5(data_out_5),
	.data_out_6(data_out_6),
	.data_out_7(data_out_7),
	.data_out_8(data_out_8),
	.data_out_9(data_out_9),
	.data_out_10(data_out_10),
	.data_out_11(data_out_11),
	.data_out_12(data_out_12),
	.data_out_13(data_out_13),
	.data_out_14(data_out_14),
	.data_out_15(data_out_15),
	.data_out_16(data_out_16),
	.data_out_17(data_out_17),
	.data_out_18(data_out_18),
	.data_out_19(data_out_19),
	.data_out_20(data_out_20),
	.data_out_21(data_out_21),
	.data_out_22(data_out_22),
	.data_out_23(data_out_23),
	.ram_block1a96(\ux0120|altsyncram_component0|auto_generated|ram_block1a96~portadataout ),
	.ram_block1a120(\ux0120|altsyncram_component0|auto_generated|ram_block1a120~portadataout ),
	.ram_block1a144(\ux0120|altsyncram_component0|auto_generated|ram_block1a144~portadataout ),
	.ram_block1a168(\ux0120|altsyncram_component0|auto_generated|ram_block1a168~portadataout ),
	.ram_block1a48(\ux0120|altsyncram_component0|auto_generated|ram_block1a48~portadataout ),
	.ram_block1a72(\ux0120|altsyncram_component0|auto_generated|ram_block1a72~portadataout ),
	.ram_block1a0(\ux0120|altsyncram_component0|auto_generated|ram_block1a0~portadataout ),
	.ram_block1a24(\ux0120|altsyncram_component0|auto_generated|ram_block1a24~portadataout ),
	.ram_block1a97(\ux0120|altsyncram_component0|auto_generated|ram_block1a97~portadataout ),
	.ram_block1a121(\ux0120|altsyncram_component0|auto_generated|ram_block1a121~portadataout ),
	.ram_block1a145(\ux0120|altsyncram_component0|auto_generated|ram_block1a145~portadataout ),
	.ram_block1a169(\ux0120|altsyncram_component0|auto_generated|ram_block1a169~portadataout ),
	.ram_block1a49(\ux0120|altsyncram_component0|auto_generated|ram_block1a49~portadataout ),
	.ram_block1a73(\ux0120|altsyncram_component0|auto_generated|ram_block1a73~portadataout ),
	.ram_block1a1(\ux0120|altsyncram_component0|auto_generated|ram_block1a1~portadataout ),
	.ram_block1a25(\ux0120|altsyncram_component0|auto_generated|ram_block1a25~portadataout ),
	.ram_block1a98(\ux0120|altsyncram_component0|auto_generated|ram_block1a98~portadataout ),
	.ram_block1a122(\ux0120|altsyncram_component0|auto_generated|ram_block1a122~portadataout ),
	.ram_block1a146(\ux0120|altsyncram_component0|auto_generated|ram_block1a146~portadataout ),
	.ram_block1a170(\ux0120|altsyncram_component0|auto_generated|ram_block1a170~portadataout ),
	.ram_block1a50(\ux0120|altsyncram_component0|auto_generated|ram_block1a50~portadataout ),
	.ram_block1a74(\ux0120|altsyncram_component0|auto_generated|ram_block1a74~portadataout ),
	.ram_block1a2(\ux0120|altsyncram_component0|auto_generated|ram_block1a2~portadataout ),
	.ram_block1a26(\ux0120|altsyncram_component0|auto_generated|ram_block1a26~portadataout ),
	.ram_block1a99(\ux0120|altsyncram_component0|auto_generated|ram_block1a99~portadataout ),
	.ram_block1a123(\ux0120|altsyncram_component0|auto_generated|ram_block1a123~portadataout ),
	.ram_block1a147(\ux0120|altsyncram_component0|auto_generated|ram_block1a147~portadataout ),
	.ram_block1a171(\ux0120|altsyncram_component0|auto_generated|ram_block1a171~portadataout ),
	.ram_block1a51(\ux0120|altsyncram_component0|auto_generated|ram_block1a51~portadataout ),
	.ram_block1a75(\ux0120|altsyncram_component0|auto_generated|ram_block1a75~portadataout ),
	.ram_block1a3(\ux0120|altsyncram_component0|auto_generated|ram_block1a3~portadataout ),
	.ram_block1a27(\ux0120|altsyncram_component0|auto_generated|ram_block1a27~portadataout ),
	.ram_block1a100(\ux0120|altsyncram_component0|auto_generated|ram_block1a100~portadataout ),
	.ram_block1a124(\ux0120|altsyncram_component0|auto_generated|ram_block1a124~portadataout ),
	.ram_block1a148(\ux0120|altsyncram_component0|auto_generated|ram_block1a148~portadataout ),
	.ram_block1a172(\ux0120|altsyncram_component0|auto_generated|ram_block1a172~portadataout ),
	.ram_block1a52(\ux0120|altsyncram_component0|auto_generated|ram_block1a52~portadataout ),
	.ram_block1a76(\ux0120|altsyncram_component0|auto_generated|ram_block1a76~portadataout ),
	.ram_block1a4(\ux0120|altsyncram_component0|auto_generated|ram_block1a4~portadataout ),
	.ram_block1a28(\ux0120|altsyncram_component0|auto_generated|ram_block1a28~portadataout ),
	.ram_block1a101(\ux0120|altsyncram_component0|auto_generated|ram_block1a101~portadataout ),
	.ram_block1a125(\ux0120|altsyncram_component0|auto_generated|ram_block1a125~portadataout ),
	.ram_block1a149(\ux0120|altsyncram_component0|auto_generated|ram_block1a149~portadataout ),
	.ram_block1a173(\ux0120|altsyncram_component0|auto_generated|ram_block1a173~portadataout ),
	.ram_block1a53(\ux0120|altsyncram_component0|auto_generated|ram_block1a53~portadataout ),
	.ram_block1a77(\ux0120|altsyncram_component0|auto_generated|ram_block1a77~portadataout ),
	.ram_block1a5(\ux0120|altsyncram_component0|auto_generated|ram_block1a5~portadataout ),
	.ram_block1a29(\ux0120|altsyncram_component0|auto_generated|ram_block1a29~portadataout ),
	.ram_block1a102(\ux0120|altsyncram_component0|auto_generated|ram_block1a102~portadataout ),
	.ram_block1a126(\ux0120|altsyncram_component0|auto_generated|ram_block1a126~portadataout ),
	.ram_block1a150(\ux0120|altsyncram_component0|auto_generated|ram_block1a150~portadataout ),
	.ram_block1a174(\ux0120|altsyncram_component0|auto_generated|ram_block1a174~portadataout ),
	.ram_block1a54(\ux0120|altsyncram_component0|auto_generated|ram_block1a54~portadataout ),
	.ram_block1a78(\ux0120|altsyncram_component0|auto_generated|ram_block1a78~portadataout ),
	.ram_block1a6(\ux0120|altsyncram_component0|auto_generated|ram_block1a6~portadataout ),
	.ram_block1a30(\ux0120|altsyncram_component0|auto_generated|ram_block1a30~portadataout ),
	.ram_block1a103(\ux0120|altsyncram_component0|auto_generated|ram_block1a103~portadataout ),
	.ram_block1a127(\ux0120|altsyncram_component0|auto_generated|ram_block1a127~portadataout ),
	.ram_block1a151(\ux0120|altsyncram_component0|auto_generated|ram_block1a151~portadataout ),
	.ram_block1a175(\ux0120|altsyncram_component0|auto_generated|ram_block1a175~portadataout ),
	.ram_block1a55(\ux0120|altsyncram_component0|auto_generated|ram_block1a55~portadataout ),
	.ram_block1a79(\ux0120|altsyncram_component0|auto_generated|ram_block1a79~portadataout ),
	.ram_block1a7(\ux0120|altsyncram_component0|auto_generated|ram_block1a7~portadataout ),
	.ram_block1a31(\ux0120|altsyncram_component0|auto_generated|ram_block1a31~portadataout ),
	.ram_block1a104(\ux0120|altsyncram_component0|auto_generated|ram_block1a104~portadataout ),
	.ram_block1a128(\ux0120|altsyncram_component0|auto_generated|ram_block1a128~portadataout ),
	.ram_block1a152(\ux0120|altsyncram_component0|auto_generated|ram_block1a152~portadataout ),
	.ram_block1a176(\ux0120|altsyncram_component0|auto_generated|ram_block1a176~portadataout ),
	.ram_block1a56(\ux0120|altsyncram_component0|auto_generated|ram_block1a56~portadataout ),
	.ram_block1a80(\ux0120|altsyncram_component0|auto_generated|ram_block1a80~portadataout ),
	.ram_block1a8(\ux0120|altsyncram_component0|auto_generated|ram_block1a8~portadataout ),
	.ram_block1a32(\ux0120|altsyncram_component0|auto_generated|ram_block1a32~portadataout ),
	.ram_block1a105(\ux0120|altsyncram_component0|auto_generated|ram_block1a105~portadataout ),
	.ram_block1a129(\ux0120|altsyncram_component0|auto_generated|ram_block1a129~portadataout ),
	.ram_block1a153(\ux0120|altsyncram_component0|auto_generated|ram_block1a153~portadataout ),
	.ram_block1a177(\ux0120|altsyncram_component0|auto_generated|ram_block1a177~portadataout ),
	.ram_block1a57(\ux0120|altsyncram_component0|auto_generated|ram_block1a57~portadataout ),
	.ram_block1a81(\ux0120|altsyncram_component0|auto_generated|ram_block1a81~portadataout ),
	.ram_block1a9(\ux0120|altsyncram_component0|auto_generated|ram_block1a9~portadataout ),
	.ram_block1a33(\ux0120|altsyncram_component0|auto_generated|ram_block1a33~portadataout ),
	.ram_block1a106(\ux0120|altsyncram_component0|auto_generated|ram_block1a106~portadataout ),
	.ram_block1a130(\ux0120|altsyncram_component0|auto_generated|ram_block1a130~portadataout ),
	.ram_block1a154(\ux0120|altsyncram_component0|auto_generated|ram_block1a154~portadataout ),
	.ram_block1a178(\ux0120|altsyncram_component0|auto_generated|ram_block1a178~portadataout ),
	.ram_block1a58(\ux0120|altsyncram_component0|auto_generated|ram_block1a58~portadataout ),
	.ram_block1a82(\ux0120|altsyncram_component0|auto_generated|ram_block1a82~portadataout ),
	.ram_block1a10(\ux0120|altsyncram_component0|auto_generated|ram_block1a10~portadataout ),
	.ram_block1a34(\ux0120|altsyncram_component0|auto_generated|ram_block1a34~portadataout ),
	.ram_block1a107(\ux0120|altsyncram_component0|auto_generated|ram_block1a107~portadataout ),
	.ram_block1a131(\ux0120|altsyncram_component0|auto_generated|ram_block1a131~portadataout ),
	.ram_block1a155(\ux0120|altsyncram_component0|auto_generated|ram_block1a155~portadataout ),
	.ram_block1a179(\ux0120|altsyncram_component0|auto_generated|ram_block1a179~portadataout ),
	.ram_block1a59(\ux0120|altsyncram_component0|auto_generated|ram_block1a59~portadataout ),
	.ram_block1a83(\ux0120|altsyncram_component0|auto_generated|ram_block1a83~portadataout ),
	.ram_block1a11(\ux0120|altsyncram_component0|auto_generated|ram_block1a11~portadataout ),
	.ram_block1a35(\ux0120|altsyncram_component0|auto_generated|ram_block1a35~portadataout ),
	.ram_block1a108(\ux0120|altsyncram_component0|auto_generated|ram_block1a108~portadataout ),
	.ram_block1a132(\ux0120|altsyncram_component0|auto_generated|ram_block1a132~portadataout ),
	.ram_block1a156(\ux0120|altsyncram_component0|auto_generated|ram_block1a156~portadataout ),
	.ram_block1a180(\ux0120|altsyncram_component0|auto_generated|ram_block1a180~portadataout ),
	.ram_block1a60(\ux0120|altsyncram_component0|auto_generated|ram_block1a60~portadataout ),
	.ram_block1a84(\ux0120|altsyncram_component0|auto_generated|ram_block1a84~portadataout ),
	.ram_block1a12(\ux0120|altsyncram_component0|auto_generated|ram_block1a12~portadataout ),
	.ram_block1a36(\ux0120|altsyncram_component0|auto_generated|ram_block1a36~portadataout ),
	.ram_block1a109(\ux0120|altsyncram_component0|auto_generated|ram_block1a109~portadataout ),
	.ram_block1a133(\ux0120|altsyncram_component0|auto_generated|ram_block1a133~portadataout ),
	.ram_block1a157(\ux0120|altsyncram_component0|auto_generated|ram_block1a157~portadataout ),
	.ram_block1a181(\ux0120|altsyncram_component0|auto_generated|ram_block1a181~portadataout ),
	.ram_block1a61(\ux0120|altsyncram_component0|auto_generated|ram_block1a61~portadataout ),
	.ram_block1a85(\ux0120|altsyncram_component0|auto_generated|ram_block1a85~portadataout ),
	.ram_block1a13(\ux0120|altsyncram_component0|auto_generated|ram_block1a13~portadataout ),
	.ram_block1a37(\ux0120|altsyncram_component0|auto_generated|ram_block1a37~portadataout ),
	.ram_block1a110(\ux0120|altsyncram_component0|auto_generated|ram_block1a110~portadataout ),
	.ram_block1a134(\ux0120|altsyncram_component0|auto_generated|ram_block1a134~portadataout ),
	.ram_block1a158(\ux0120|altsyncram_component0|auto_generated|ram_block1a158~portadataout ),
	.ram_block1a182(\ux0120|altsyncram_component0|auto_generated|ram_block1a182~portadataout ),
	.ram_block1a62(\ux0120|altsyncram_component0|auto_generated|ram_block1a62~portadataout ),
	.ram_block1a86(\ux0120|altsyncram_component0|auto_generated|ram_block1a86~portadataout ),
	.ram_block1a14(\ux0120|altsyncram_component0|auto_generated|ram_block1a14~portadataout ),
	.ram_block1a38(\ux0120|altsyncram_component0|auto_generated|ram_block1a38~portadataout ),
	.ram_block1a111(\ux0120|altsyncram_component0|auto_generated|ram_block1a111~portadataout ),
	.ram_block1a135(\ux0120|altsyncram_component0|auto_generated|ram_block1a135~portadataout ),
	.ram_block1a159(\ux0120|altsyncram_component0|auto_generated|ram_block1a159~portadataout ),
	.ram_block1a183(\ux0120|altsyncram_component0|auto_generated|ram_block1a183~portadataout ),
	.ram_block1a63(\ux0120|altsyncram_component0|auto_generated|ram_block1a63~portadataout ),
	.ram_block1a87(\ux0120|altsyncram_component0|auto_generated|ram_block1a87~portadataout ),
	.ram_block1a15(\ux0120|altsyncram_component0|auto_generated|ram_block1a15~portadataout ),
	.ram_block1a39(\ux0120|altsyncram_component0|auto_generated|ram_block1a39~portadataout ),
	.ram_block1a112(\ux0120|altsyncram_component0|auto_generated|ram_block1a112~portadataout ),
	.ram_block1a136(\ux0120|altsyncram_component0|auto_generated|ram_block1a136~portadataout ),
	.ram_block1a160(\ux0120|altsyncram_component0|auto_generated|ram_block1a160~portadataout ),
	.ram_block1a184(\ux0120|altsyncram_component0|auto_generated|ram_block1a184~portadataout ),
	.ram_block1a64(\ux0120|altsyncram_component0|auto_generated|ram_block1a64~portadataout ),
	.ram_block1a88(\ux0120|altsyncram_component0|auto_generated|ram_block1a88~portadataout ),
	.ram_block1a16(\ux0120|altsyncram_component0|auto_generated|ram_block1a16~portadataout ),
	.ram_block1a40(\ux0120|altsyncram_component0|auto_generated|ram_block1a40~portadataout ),
	.ram_block1a113(\ux0120|altsyncram_component0|auto_generated|ram_block1a113~portadataout ),
	.ram_block1a137(\ux0120|altsyncram_component0|auto_generated|ram_block1a137~portadataout ),
	.ram_block1a161(\ux0120|altsyncram_component0|auto_generated|ram_block1a161~portadataout ),
	.ram_block1a185(\ux0120|altsyncram_component0|auto_generated|ram_block1a185~portadataout ),
	.ram_block1a65(\ux0120|altsyncram_component0|auto_generated|ram_block1a65~portadataout ),
	.ram_block1a89(\ux0120|altsyncram_component0|auto_generated|ram_block1a89~portadataout ),
	.ram_block1a17(\ux0120|altsyncram_component0|auto_generated|ram_block1a17~portadataout ),
	.ram_block1a41(\ux0120|altsyncram_component0|auto_generated|ram_block1a41~portadataout ),
	.ram_block1a114(\ux0120|altsyncram_component0|auto_generated|ram_block1a114~portadataout ),
	.ram_block1a138(\ux0120|altsyncram_component0|auto_generated|ram_block1a138~portadataout ),
	.ram_block1a162(\ux0120|altsyncram_component0|auto_generated|ram_block1a162~portadataout ),
	.ram_block1a186(\ux0120|altsyncram_component0|auto_generated|ram_block1a186~portadataout ),
	.ram_block1a66(\ux0120|altsyncram_component0|auto_generated|ram_block1a66~portadataout ),
	.ram_block1a90(\ux0120|altsyncram_component0|auto_generated|ram_block1a90~portadataout ),
	.ram_block1a18(\ux0120|altsyncram_component0|auto_generated|ram_block1a18~portadataout ),
	.ram_block1a42(\ux0120|altsyncram_component0|auto_generated|ram_block1a42~portadataout ),
	.ram_block1a115(\ux0120|altsyncram_component0|auto_generated|ram_block1a115~portadataout ),
	.ram_block1a139(\ux0120|altsyncram_component0|auto_generated|ram_block1a139~portadataout ),
	.ram_block1a163(\ux0120|altsyncram_component0|auto_generated|ram_block1a163~portadataout ),
	.ram_block1a187(\ux0120|altsyncram_component0|auto_generated|ram_block1a187~portadataout ),
	.ram_block1a67(\ux0120|altsyncram_component0|auto_generated|ram_block1a67~portadataout ),
	.ram_block1a91(\ux0120|altsyncram_component0|auto_generated|ram_block1a91~portadataout ),
	.ram_block1a19(\ux0120|altsyncram_component0|auto_generated|ram_block1a19~portadataout ),
	.ram_block1a43(\ux0120|altsyncram_component0|auto_generated|ram_block1a43~portadataout ),
	.ram_block1a116(\ux0120|altsyncram_component0|auto_generated|ram_block1a116~portadataout ),
	.ram_block1a140(\ux0120|altsyncram_component0|auto_generated|ram_block1a140~portadataout ),
	.ram_block1a164(\ux0120|altsyncram_component0|auto_generated|ram_block1a164~portadataout ),
	.ram_block1a188(\ux0120|altsyncram_component0|auto_generated|ram_block1a188~portadataout ),
	.ram_block1a68(\ux0120|altsyncram_component0|auto_generated|ram_block1a68~portadataout ),
	.ram_block1a92(\ux0120|altsyncram_component0|auto_generated|ram_block1a92~portadataout ),
	.ram_block1a20(\ux0120|altsyncram_component0|auto_generated|ram_block1a20~portadataout ),
	.ram_block1a44(\ux0120|altsyncram_component0|auto_generated|ram_block1a44~portadataout ),
	.ram_block1a117(\ux0120|altsyncram_component0|auto_generated|ram_block1a117~portadataout ),
	.ram_block1a141(\ux0120|altsyncram_component0|auto_generated|ram_block1a141~portadataout ),
	.ram_block1a165(\ux0120|altsyncram_component0|auto_generated|ram_block1a165~portadataout ),
	.ram_block1a189(\ux0120|altsyncram_component0|auto_generated|ram_block1a189~portadataout ),
	.ram_block1a69(\ux0120|altsyncram_component0|auto_generated|ram_block1a69~portadataout ),
	.ram_block1a93(\ux0120|altsyncram_component0|auto_generated|ram_block1a93~portadataout ),
	.ram_block1a21(\ux0120|altsyncram_component0|auto_generated|ram_block1a21~portadataout ),
	.ram_block1a45(\ux0120|altsyncram_component0|auto_generated|ram_block1a45~portadataout ),
	.ram_block1a118(\ux0120|altsyncram_component0|auto_generated|ram_block1a118~portadataout ),
	.ram_block1a142(\ux0120|altsyncram_component0|auto_generated|ram_block1a142~portadataout ),
	.ram_block1a166(\ux0120|altsyncram_component0|auto_generated|ram_block1a166~portadataout ),
	.ram_block1a190(\ux0120|altsyncram_component0|auto_generated|ram_block1a190~portadataout ),
	.ram_block1a70(\ux0120|altsyncram_component0|auto_generated|ram_block1a70~portadataout ),
	.ram_block1a94(\ux0120|altsyncram_component0|auto_generated|ram_block1a94~portadataout ),
	.ram_block1a22(\ux0120|altsyncram_component0|auto_generated|ram_block1a22~portadataout ),
	.ram_block1a46(\ux0120|altsyncram_component0|auto_generated|ram_block1a46~portadataout ),
	.ram_block1a119(\ux0120|altsyncram_component0|auto_generated|ram_block1a119~portadataout ),
	.ram_block1a143(\ux0120|altsyncram_component0|auto_generated|ram_block1a143~portadataout ),
	.ram_block1a167(\ux0120|altsyncram_component0|auto_generated|ram_block1a167~portadataout ),
	.ram_block1a191(\ux0120|altsyncram_component0|auto_generated|ram_block1a191~portadataout ),
	.ram_block1a71(\ux0120|altsyncram_component0|auto_generated|ram_block1a71~portadataout ),
	.ram_block1a95(\ux0120|altsyncram_component0|auto_generated|ram_block1a95~portadataout ),
	.ram_block1a23(\ux0120|altsyncram_component0|auto_generated|ram_block1a23~portadataout ),
	.ram_block1a47(\ux0120|altsyncram_component0|auto_generated|ram_block1a47~portadataout ),
	.out_address_reg_a_2(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[2]~q ),
	.out_address_reg_a_0(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[0]~q ),
	.out_address_reg_a_1(\ux0120|altsyncram_component0|auto_generated|out_address_reg_a[1]~q ),
	.data_out_121(\ux122|data_out[12]~3_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module sine_asj_altqmcpipe (
	data_out_12,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_31,
	pipeline_dffe_15,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_14,
	pipeline_dffe_161,
	pipeline_dffe_13,
	pipeline_dffe_171,
	pipeline_dffe_181,
	pipeline_dffe_191,
	pipeline_dffe_201,
	pipeline_dffe_211,
	pipeline_dffe_221,
	pipeline_dffe_231,
	pipeline_dffe_241,
	pipeline_dffe_251,
	pipeline_dffe_261,
	pipeline_dffe_271,
	pipeline_dffe_281,
	pipeline_dffe_311,
	pipeline_dffe_151,
	pipeline_dffe_12,
	pipeline_dffe_291,
	pipeline_dffe_301,
	pipeline_dffe_141,
	pipeline_dffe_11,
	pipeline_dffe_131,
	pipeline_dffe_121,
	pipeline_dffe_111,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	data_out_12;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_31;
output 	pipeline_dffe_15;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_14;
input 	pipeline_dffe_161;
output 	pipeline_dffe_13;
input 	pipeline_dffe_171;
input 	pipeline_dffe_181;
input 	pipeline_dffe_191;
input 	pipeline_dffe_201;
input 	pipeline_dffe_211;
input 	pipeline_dffe_221;
input 	pipeline_dffe_231;
input 	pipeline_dffe_241;
input 	pipeline_dffe_251;
input 	pipeline_dffe_261;
input 	pipeline_dffe_271;
input 	pipeline_dffe_281;
input 	pipeline_dffe_311;
input 	pipeline_dffe_151;
output 	pipeline_dffe_12;
input 	pipeline_dffe_291;
input 	pipeline_dffe_301;
input 	pipeline_dffe_141;
output 	pipeline_dffe_11;
input 	pipeline_dffe_131;
input 	pipeline_dffe_121;
input 	pipeline_dffe_111;
input 	pipeline_dffe_10;
input 	pipeline_dffe_9;
input 	pipeline_dffe_8;
input 	pipeline_dffe_7;
input 	pipeline_dffe_6;
input 	pipeline_dffe_5;
input 	pipeline_dffe_4;
input 	pipeline_dffe_3;
input 	pipeline_dffe_2;
input 	pipeline_dffe_1;
input 	pipeline_dffe_0;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \phi_int_arr_reg[16]~q ;
wire \phi_int_arr_reg[17]~q ;
wire \phi_int_arr_reg[18]~q ;
wire \phi_int_arr_reg[19]~q ;
wire \phi_int_arr_reg[20]~q ;
wire \phi_int_arr_reg[21]~q ;
wire \phi_int_arr_reg[22]~q ;
wire \phi_int_arr_reg[23]~q ;
wire \phi_int_arr_reg[24]~q ;
wire \phi_int_arr_reg[25]~q ;
wire \phi_int_arr_reg[26]~q ;
wire \phi_int_arr_reg[27]~q ;
wire \phi_int_arr_reg[28]~q ;
wire \phi_int_arr_reg[31]~q ;
wire \phi_int_arr_reg[15]~q ;
wire \phi_int_arr_reg[29]~q ;
wire \phi_int_arr_reg[30]~q ;
wire \phi_int_arr_reg[14]~q ;
wire \phi_int_arr_reg[13]~q ;
wire \phi_int_arr_reg[12]~q ;
wire \phi_int_arr_reg[11]~q ;
wire \phi_int_arr_reg[10]~q ;
wire \phi_int_arr_reg[9]~q ;
wire \phi_int_arr_reg[8]~q ;
wire \phi_int_arr_reg[7]~q ;
wire \phi_int_arr_reg[6]~q ;
wire \phi_int_arr_reg[5]~q ;
wire \phi_int_arr_reg[4]~q ;
wire \phi_int_arr_reg[3]~q ;
wire \phi_int_arr_reg[2]~q ;
wire \phi_int_arr_reg[1]~q ;
wire \phi_int_arr_reg[0]~q ;


sine_lpm_add_sub_1 acc(
	.phi_int_arr_reg_16(\phi_int_arr_reg[16]~q ),
	.phi_int_arr_reg_17(\phi_int_arr_reg[17]~q ),
	.phi_int_arr_reg_18(\phi_int_arr_reg[18]~q ),
	.phi_int_arr_reg_19(\phi_int_arr_reg[19]~q ),
	.phi_int_arr_reg_20(\phi_int_arr_reg[20]~q ),
	.phi_int_arr_reg_21(\phi_int_arr_reg[21]~q ),
	.phi_int_arr_reg_22(\phi_int_arr_reg[22]~q ),
	.phi_int_arr_reg_23(\phi_int_arr_reg[23]~q ),
	.phi_int_arr_reg_24(\phi_int_arr_reg[24]~q ),
	.phi_int_arr_reg_25(\phi_int_arr_reg[25]~q ),
	.phi_int_arr_reg_26(\phi_int_arr_reg[26]~q ),
	.phi_int_arr_reg_27(\phi_int_arr_reg[27]~q ),
	.phi_int_arr_reg_28(\phi_int_arr_reg[28]~q ),
	.phi_int_arr_reg_31(\phi_int_arr_reg[31]~q ),
	.phi_int_arr_reg_15(\phi_int_arr_reg[15]~q ),
	.phi_int_arr_reg_29(\phi_int_arr_reg[29]~q ),
	.phi_int_arr_reg_30(\phi_int_arr_reg[30]~q ),
	.phi_int_arr_reg_14(\phi_int_arr_reg[14]~q ),
	.phi_int_arr_reg_13(\phi_int_arr_reg[13]~q ),
	.phi_int_arr_reg_12(\phi_int_arr_reg[12]~q ),
	.phi_int_arr_reg_11(\phi_int_arr_reg[11]~q ),
	.phi_int_arr_reg_10(\phi_int_arr_reg[10]~q ),
	.phi_int_arr_reg_9(\phi_int_arr_reg[9]~q ),
	.phi_int_arr_reg_8(\phi_int_arr_reg[8]~q ),
	.phi_int_arr_reg_7(\phi_int_arr_reg[7]~q ),
	.phi_int_arr_reg_6(\phi_int_arr_reg[6]~q ),
	.phi_int_arr_reg_5(\phi_int_arr_reg[5]~q ),
	.phi_int_arr_reg_4(\phi_int_arr_reg[4]~q ),
	.phi_int_arr_reg_3(\phi_int_arr_reg[3]~q ),
	.phi_int_arr_reg_2(\phi_int_arr_reg[2]~q ),
	.phi_int_arr_reg_1(\phi_int_arr_reg[1]~q ),
	.phi_int_arr_reg_0(\phi_int_arr_reg[0]~q ),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \phi_int_arr_reg[16] (
	.clk(clk),
	.d(pipeline_dffe_161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[16]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[16] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[16] .power_up = "low";

dffeas \phi_int_arr_reg[17] (
	.clk(clk),
	.d(pipeline_dffe_171),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[17]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[17] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[17] .power_up = "low";

dffeas \phi_int_arr_reg[18] (
	.clk(clk),
	.d(pipeline_dffe_181),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[18]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[18] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[18] .power_up = "low";

dffeas \phi_int_arr_reg[19] (
	.clk(clk),
	.d(pipeline_dffe_191),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[19]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[19] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[19] .power_up = "low";

dffeas \phi_int_arr_reg[20] (
	.clk(clk),
	.d(pipeline_dffe_201),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[20]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[20] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[20] .power_up = "low";

dffeas \phi_int_arr_reg[21] (
	.clk(clk),
	.d(pipeline_dffe_211),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[21]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[21] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[21] .power_up = "low";

dffeas \phi_int_arr_reg[22] (
	.clk(clk),
	.d(pipeline_dffe_221),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[22]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[22] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[22] .power_up = "low";

dffeas \phi_int_arr_reg[23] (
	.clk(clk),
	.d(pipeline_dffe_231),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[23]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[23] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[23] .power_up = "low";

dffeas \phi_int_arr_reg[24] (
	.clk(clk),
	.d(pipeline_dffe_241),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[24]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[24] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[24] .power_up = "low";

dffeas \phi_int_arr_reg[25] (
	.clk(clk),
	.d(pipeline_dffe_251),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[25]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[25] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[25] .power_up = "low";

dffeas \phi_int_arr_reg[26] (
	.clk(clk),
	.d(pipeline_dffe_261),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[26]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[26] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[26] .power_up = "low";

dffeas \phi_int_arr_reg[27] (
	.clk(clk),
	.d(pipeline_dffe_271),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[27]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[27] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[27] .power_up = "low";

dffeas \phi_int_arr_reg[28] (
	.clk(clk),
	.d(pipeline_dffe_281),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[28]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[28] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[28] .power_up = "low";

dffeas \phi_int_arr_reg[31] (
	.clk(clk),
	.d(pipeline_dffe_311),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[31]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[31] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[31] .power_up = "low";

dffeas \phi_int_arr_reg[15] (
	.clk(clk),
	.d(pipeline_dffe_151),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[15]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[15] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[15] .power_up = "low";

dffeas \phi_int_arr_reg[29] (
	.clk(clk),
	.d(pipeline_dffe_291),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[29]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[29] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[29] .power_up = "low";

dffeas \phi_int_arr_reg[30] (
	.clk(clk),
	.d(pipeline_dffe_301),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[30]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[30] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[30] .power_up = "low";

dffeas \phi_int_arr_reg[14] (
	.clk(clk),
	.d(pipeline_dffe_141),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[14]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[14] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[14] .power_up = "low";

dffeas \phi_int_arr_reg[13] (
	.clk(clk),
	.d(pipeline_dffe_131),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[13]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[13] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[13] .power_up = "low";

dffeas \phi_int_arr_reg[12] (
	.clk(clk),
	.d(pipeline_dffe_121),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[12]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[12] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[12] .power_up = "low";

dffeas \phi_int_arr_reg[11] (
	.clk(clk),
	.d(pipeline_dffe_111),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[11]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[11] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[11] .power_up = "low";

dffeas \phi_int_arr_reg[10] (
	.clk(clk),
	.d(pipeline_dffe_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[10]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[10] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[10] .power_up = "low";

dffeas \phi_int_arr_reg[9] (
	.clk(clk),
	.d(pipeline_dffe_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[9]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[9] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[9] .power_up = "low";

dffeas \phi_int_arr_reg[8] (
	.clk(clk),
	.d(pipeline_dffe_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[8]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[8] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[8] .power_up = "low";

dffeas \phi_int_arr_reg[7] (
	.clk(clk),
	.d(pipeline_dffe_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[7]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[7] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[7] .power_up = "low";

dffeas \phi_int_arr_reg[6] (
	.clk(clk),
	.d(pipeline_dffe_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[6]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[6] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[6] .power_up = "low";

dffeas \phi_int_arr_reg[5] (
	.clk(clk),
	.d(pipeline_dffe_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[5]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[5] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[5] .power_up = "low";

dffeas \phi_int_arr_reg[4] (
	.clk(clk),
	.d(pipeline_dffe_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[4]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[4] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[4] .power_up = "low";

dffeas \phi_int_arr_reg[3] (
	.clk(clk),
	.d(pipeline_dffe_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[3]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[3] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[3] .power_up = "low";

dffeas \phi_int_arr_reg[2] (
	.clk(clk),
	.d(pipeline_dffe_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[2]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[2] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[2] .power_up = "low";

dffeas \phi_int_arr_reg[1] (
	.clk(clk),
	.d(pipeline_dffe_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[1]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[1] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[1] .power_up = "low";

dffeas \phi_int_arr_reg[0] (
	.clk(clk),
	.d(pipeline_dffe_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_int_arr_reg[0]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[0] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[0] .power_up = "low";

endmodule

module sine_lpm_add_sub_1 (
	phi_int_arr_reg_16,
	phi_int_arr_reg_17,
	phi_int_arr_reg_18,
	phi_int_arr_reg_19,
	phi_int_arr_reg_20,
	phi_int_arr_reg_21,
	phi_int_arr_reg_22,
	phi_int_arr_reg_23,
	phi_int_arr_reg_24,
	phi_int_arr_reg_25,
	phi_int_arr_reg_26,
	phi_int_arr_reg_27,
	phi_int_arr_reg_28,
	phi_int_arr_reg_31,
	phi_int_arr_reg_15,
	phi_int_arr_reg_29,
	phi_int_arr_reg_30,
	phi_int_arr_reg_14,
	phi_int_arr_reg_13,
	phi_int_arr_reg_12,
	phi_int_arr_reg_11,
	phi_int_arr_reg_10,
	phi_int_arr_reg_9,
	phi_int_arr_reg_8,
	phi_int_arr_reg_7,
	phi_int_arr_reg_6,
	phi_int_arr_reg_5,
	phi_int_arr_reg_4,
	phi_int_arr_reg_3,
	phi_int_arr_reg_2,
	phi_int_arr_reg_1,
	phi_int_arr_reg_0,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_31,
	pipeline_dffe_15,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	phi_int_arr_reg_16;
input 	phi_int_arr_reg_17;
input 	phi_int_arr_reg_18;
input 	phi_int_arr_reg_19;
input 	phi_int_arr_reg_20;
input 	phi_int_arr_reg_21;
input 	phi_int_arr_reg_22;
input 	phi_int_arr_reg_23;
input 	phi_int_arr_reg_24;
input 	phi_int_arr_reg_25;
input 	phi_int_arr_reg_26;
input 	phi_int_arr_reg_27;
input 	phi_int_arr_reg_28;
input 	phi_int_arr_reg_31;
input 	phi_int_arr_reg_15;
input 	phi_int_arr_reg_29;
input 	phi_int_arr_reg_30;
input 	phi_int_arr_reg_14;
input 	phi_int_arr_reg_13;
input 	phi_int_arr_reg_12;
input 	phi_int_arr_reg_11;
input 	phi_int_arr_reg_10;
input 	phi_int_arr_reg_9;
input 	phi_int_arr_reg_8;
input 	phi_int_arr_reg_7;
input 	phi_int_arr_reg_6;
input 	phi_int_arr_reg_5;
input 	phi_int_arr_reg_4;
input 	phi_int_arr_reg_3;
input 	phi_int_arr_reg_2;
input 	phi_int_arr_reg_1;
input 	phi_int_arr_reg_0;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_31;
output 	pipeline_dffe_15;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_add_sub_hth auto_generated(
	.phi_int_arr_reg_16(phi_int_arr_reg_16),
	.phi_int_arr_reg_17(phi_int_arr_reg_17),
	.phi_int_arr_reg_18(phi_int_arr_reg_18),
	.phi_int_arr_reg_19(phi_int_arr_reg_19),
	.phi_int_arr_reg_20(phi_int_arr_reg_20),
	.phi_int_arr_reg_21(phi_int_arr_reg_21),
	.phi_int_arr_reg_22(phi_int_arr_reg_22),
	.phi_int_arr_reg_23(phi_int_arr_reg_23),
	.phi_int_arr_reg_24(phi_int_arr_reg_24),
	.phi_int_arr_reg_25(phi_int_arr_reg_25),
	.phi_int_arr_reg_26(phi_int_arr_reg_26),
	.phi_int_arr_reg_27(phi_int_arr_reg_27),
	.phi_int_arr_reg_28(phi_int_arr_reg_28),
	.phi_int_arr_reg_31(phi_int_arr_reg_31),
	.phi_int_arr_reg_15(phi_int_arr_reg_15),
	.phi_int_arr_reg_29(phi_int_arr_reg_29),
	.phi_int_arr_reg_30(phi_int_arr_reg_30),
	.phi_int_arr_reg_14(phi_int_arr_reg_14),
	.phi_int_arr_reg_13(phi_int_arr_reg_13),
	.phi_int_arr_reg_12(phi_int_arr_reg_12),
	.phi_int_arr_reg_11(phi_int_arr_reg_11),
	.phi_int_arr_reg_10(phi_int_arr_reg_10),
	.phi_int_arr_reg_9(phi_int_arr_reg_9),
	.phi_int_arr_reg_8(phi_int_arr_reg_8),
	.phi_int_arr_reg_7(phi_int_arr_reg_7),
	.phi_int_arr_reg_6(phi_int_arr_reg_6),
	.phi_int_arr_reg_5(phi_int_arr_reg_5),
	.phi_int_arr_reg_4(phi_int_arr_reg_4),
	.phi_int_arr_reg_3(phi_int_arr_reg_3),
	.phi_int_arr_reg_2(phi_int_arr_reg_2),
	.phi_int_arr_reg_1(phi_int_arr_reg_1),
	.phi_int_arr_reg_0(phi_int_arr_reg_0),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module sine_add_sub_hth (
	phi_int_arr_reg_16,
	phi_int_arr_reg_17,
	phi_int_arr_reg_18,
	phi_int_arr_reg_19,
	phi_int_arr_reg_20,
	phi_int_arr_reg_21,
	phi_int_arr_reg_22,
	phi_int_arr_reg_23,
	phi_int_arr_reg_24,
	phi_int_arr_reg_25,
	phi_int_arr_reg_26,
	phi_int_arr_reg_27,
	phi_int_arr_reg_28,
	phi_int_arr_reg_31,
	phi_int_arr_reg_15,
	phi_int_arr_reg_29,
	phi_int_arr_reg_30,
	phi_int_arr_reg_14,
	phi_int_arr_reg_13,
	phi_int_arr_reg_12,
	phi_int_arr_reg_11,
	phi_int_arr_reg_10,
	phi_int_arr_reg_9,
	phi_int_arr_reg_8,
	phi_int_arr_reg_7,
	phi_int_arr_reg_6,
	phi_int_arr_reg_5,
	phi_int_arr_reg_4,
	phi_int_arr_reg_3,
	phi_int_arr_reg_2,
	phi_int_arr_reg_1,
	phi_int_arr_reg_0,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_31,
	pipeline_dffe_15,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	phi_int_arr_reg_16;
input 	phi_int_arr_reg_17;
input 	phi_int_arr_reg_18;
input 	phi_int_arr_reg_19;
input 	phi_int_arr_reg_20;
input 	phi_int_arr_reg_21;
input 	phi_int_arr_reg_22;
input 	phi_int_arr_reg_23;
input 	phi_int_arr_reg_24;
input 	phi_int_arr_reg_25;
input 	phi_int_arr_reg_26;
input 	phi_int_arr_reg_27;
input 	phi_int_arr_reg_28;
input 	phi_int_arr_reg_31;
input 	phi_int_arr_reg_15;
input 	phi_int_arr_reg_29;
input 	phi_int_arr_reg_30;
input 	phi_int_arr_reg_14;
input 	phi_int_arr_reg_13;
input 	phi_int_arr_reg_12;
input 	phi_int_arr_reg_11;
input 	phi_int_arr_reg_10;
input 	phi_int_arr_reg_9;
input 	phi_int_arr_reg_8;
input 	phi_int_arr_reg_7;
input 	phi_int_arr_reg_6;
input 	phi_int_arr_reg_5;
input 	phi_int_arr_reg_4;
input 	phi_int_arr_reg_3;
input 	phi_int_arr_reg_2;
input 	phi_int_arr_reg_1;
input 	phi_int_arr_reg_0;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_31;
output 	pipeline_dffe_15;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~125_sumout ;
wire \pipeline_dffe[0]~q ;
wire \op_1~126 ;
wire \op_1~121_sumout ;
wire \pipeline_dffe[1]~q ;
wire \op_1~122 ;
wire \op_1~117_sumout ;
wire \pipeline_dffe[2]~q ;
wire \op_1~118 ;
wire \op_1~113_sumout ;
wire \pipeline_dffe[3]~q ;
wire \op_1~114 ;
wire \op_1~109_sumout ;
wire \pipeline_dffe[4]~q ;
wire \op_1~110 ;
wire \op_1~105_sumout ;
wire \pipeline_dffe[5]~q ;
wire \op_1~106 ;
wire \op_1~101_sumout ;
wire \pipeline_dffe[6]~q ;
wire \op_1~102 ;
wire \op_1~97_sumout ;
wire \pipeline_dffe[7]~q ;
wire \op_1~98 ;
wire \op_1~93_sumout ;
wire \pipeline_dffe[8]~q ;
wire \op_1~94 ;
wire \op_1~89_sumout ;
wire \pipeline_dffe[9]~q ;
wire \op_1~90 ;
wire \op_1~85_sumout ;
wire \pipeline_dffe[10]~q ;
wire \op_1~86 ;
wire \op_1~82 ;
wire \op_1~78 ;
wire \op_1~74 ;
wire \op_1~70 ;
wire \op_1~58 ;
wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~6 ;
wire \op_1~9_sumout ;
wire \op_1~10 ;
wire \op_1~13_sumout ;
wire \op_1~14 ;
wire \op_1~17_sumout ;
wire \op_1~18 ;
wire \op_1~21_sumout ;
wire \op_1~22 ;
wire \op_1~25_sumout ;
wire \op_1~26 ;
wire \op_1~29_sumout ;
wire \op_1~30 ;
wire \op_1~33_sumout ;
wire \op_1~34 ;
wire \op_1~37_sumout ;
wire \op_1~38 ;
wire \op_1~41_sumout ;
wire \op_1~42 ;
wire \op_1~45_sumout ;
wire \op_1~46 ;
wire \op_1~49_sumout ;
wire \op_1~50 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~73_sumout ;
wire \op_1~77_sumout ;
wire \op_1~81_sumout ;


dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[18] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \pipeline_dffe[18] .is_wysiwyg = "true";
defparam \pipeline_dffe[18] .power_up = "low";

dffeas \pipeline_dffe[19] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \pipeline_dffe[19] .is_wysiwyg = "true";
defparam \pipeline_dffe[19] .power_up = "low";

dffeas \pipeline_dffe[20] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_20),
	.prn(vcc));
defparam \pipeline_dffe[20] .is_wysiwyg = "true";
defparam \pipeline_dffe[20] .power_up = "low";

dffeas \pipeline_dffe[21] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_21),
	.prn(vcc));
defparam \pipeline_dffe[21] .is_wysiwyg = "true";
defparam \pipeline_dffe[21] .power_up = "low";

dffeas \pipeline_dffe[22] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_22),
	.prn(vcc));
defparam \pipeline_dffe[22] .is_wysiwyg = "true";
defparam \pipeline_dffe[22] .power_up = "low";

dffeas \pipeline_dffe[23] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_23),
	.prn(vcc));
defparam \pipeline_dffe[23] .is_wysiwyg = "true";
defparam \pipeline_dffe[23] .power_up = "low";

dffeas \pipeline_dffe[24] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_24),
	.prn(vcc));
defparam \pipeline_dffe[24] .is_wysiwyg = "true";
defparam \pipeline_dffe[24] .power_up = "low";

dffeas \pipeline_dffe[25] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_25),
	.prn(vcc));
defparam \pipeline_dffe[25] .is_wysiwyg = "true";
defparam \pipeline_dffe[25] .power_up = "low";

dffeas \pipeline_dffe[26] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_26),
	.prn(vcc));
defparam \pipeline_dffe[26] .is_wysiwyg = "true";
defparam \pipeline_dffe[26] .power_up = "low";

dffeas \pipeline_dffe[27] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_27),
	.prn(vcc));
defparam \pipeline_dffe[27] .is_wysiwyg = "true";
defparam \pipeline_dffe[27] .power_up = "low";

dffeas \pipeline_dffe[28] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_28),
	.prn(vcc));
defparam \pipeline_dffe[28] .is_wysiwyg = "true";
defparam \pipeline_dffe[28] .power_up = "low";

dffeas \pipeline_dffe[31] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_31),
	.prn(vcc));
defparam \pipeline_dffe[31] .is_wysiwyg = "true";
defparam \pipeline_dffe[31] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[29] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_29),
	.prn(vcc));
defparam \pipeline_dffe[29] .is_wysiwyg = "true";
defparam \pipeline_dffe[29] .power_up = "low";

dffeas \pipeline_dffe[30] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_30),
	.prn(vcc));
defparam \pipeline_dffe[30] .is_wysiwyg = "true";
defparam \pipeline_dffe[30] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~73_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~77_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~81_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

cyclonev_lcell_comb \op_1~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_0),
	.datae(gnd),
	.dataf(!\pipeline_dffe[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~125_sumout ),
	.cout(\op_1~126 ),
	.shareout());
defparam \op_1~125 .extended_lut = "off";
defparam \op_1~125 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~125 .shared_arith = "off";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~125_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[0]~q ),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

cyclonev_lcell_comb \op_1~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_1),
	.datae(gnd),
	.dataf(!\pipeline_dffe[1]~q ),
	.datag(gnd),
	.cin(\op_1~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~121_sumout ),
	.cout(\op_1~122 ),
	.shareout());
defparam \op_1~121 .extended_lut = "off";
defparam \op_1~121 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~121 .shared_arith = "off";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~121_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[1]~q ),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

cyclonev_lcell_comb \op_1~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_2),
	.datae(gnd),
	.dataf(!\pipeline_dffe[2]~q ),
	.datag(gnd),
	.cin(\op_1~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~117_sumout ),
	.cout(\op_1~118 ),
	.shareout());
defparam \op_1~117 .extended_lut = "off";
defparam \op_1~117 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~117 .shared_arith = "off";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~117_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[2]~q ),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

cyclonev_lcell_comb \op_1~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_3),
	.datae(gnd),
	.dataf(!\pipeline_dffe[3]~q ),
	.datag(gnd),
	.cin(\op_1~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~113_sumout ),
	.cout(\op_1~114 ),
	.shareout());
defparam \op_1~113 .extended_lut = "off";
defparam \op_1~113 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~113 .shared_arith = "off";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~113_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[3]~q ),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

cyclonev_lcell_comb \op_1~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_4),
	.datae(gnd),
	.dataf(!\pipeline_dffe[4]~q ),
	.datag(gnd),
	.cin(\op_1~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~109_sumout ),
	.cout(\op_1~110 ),
	.shareout());
defparam \op_1~109 .extended_lut = "off";
defparam \op_1~109 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~109 .shared_arith = "off";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~109_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[4]~q ),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

cyclonev_lcell_comb \op_1~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_5),
	.datae(gnd),
	.dataf(!\pipeline_dffe[5]~q ),
	.datag(gnd),
	.cin(\op_1~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~105_sumout ),
	.cout(\op_1~106 ),
	.shareout());
defparam \op_1~105 .extended_lut = "off";
defparam \op_1~105 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~105 .shared_arith = "off";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~105_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[5]~q ),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

cyclonev_lcell_comb \op_1~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_6),
	.datae(gnd),
	.dataf(!\pipeline_dffe[6]~q ),
	.datag(gnd),
	.cin(\op_1~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~101_sumout ),
	.cout(\op_1~102 ),
	.shareout());
defparam \op_1~101 .extended_lut = "off";
defparam \op_1~101 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~101 .shared_arith = "off";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~101_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[6]~q ),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

cyclonev_lcell_comb \op_1~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_7),
	.datae(gnd),
	.dataf(!\pipeline_dffe[7]~q ),
	.datag(gnd),
	.cin(\op_1~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~97_sumout ),
	.cout(\op_1~98 ),
	.shareout());
defparam \op_1~97 .extended_lut = "off";
defparam \op_1~97 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~97 .shared_arith = "off";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~97_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[7]~q ),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

cyclonev_lcell_comb \op_1~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_8),
	.datae(gnd),
	.dataf(!\pipeline_dffe[8]~q ),
	.datag(gnd),
	.cin(\op_1~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~93_sumout ),
	.cout(\op_1~94 ),
	.shareout());
defparam \op_1~93 .extended_lut = "off";
defparam \op_1~93 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~93 .shared_arith = "off";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~93_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[8]~q ),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

cyclonev_lcell_comb \op_1~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_9),
	.datae(gnd),
	.dataf(!\pipeline_dffe[9]~q ),
	.datag(gnd),
	.cin(\op_1~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~89_sumout ),
	.cout(\op_1~90 ),
	.shareout());
defparam \op_1~89 .extended_lut = "off";
defparam \op_1~89 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~89 .shared_arith = "off";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~89_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[9]~q ),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

cyclonev_lcell_comb \op_1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_10),
	.datae(gnd),
	.dataf(!\pipeline_dffe[10]~q ),
	.datag(gnd),
	.cin(\op_1~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~85_sumout ),
	.cout(\op_1~86 ),
	.shareout());
defparam \op_1~85 .extended_lut = "off";
defparam \op_1~85 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~85 .shared_arith = "off";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~85_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[10]~q ),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

cyclonev_lcell_comb \op_1~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_11),
	.datae(gnd),
	.dataf(!pipeline_dffe_11),
	.datag(gnd),
	.cin(\op_1~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~81_sumout ),
	.cout(\op_1~82 ),
	.shareout());
defparam \op_1~81 .extended_lut = "off";
defparam \op_1~81 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~81 .shared_arith = "off";

cyclonev_lcell_comb \op_1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_12),
	.datae(gnd),
	.dataf(!pipeline_dffe_12),
	.datag(gnd),
	.cin(\op_1~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~77_sumout ),
	.cout(\op_1~78 ),
	.shareout());
defparam \op_1~77 .extended_lut = "off";
defparam \op_1~77 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~77 .shared_arith = "off";

cyclonev_lcell_comb \op_1~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_13),
	.datae(gnd),
	.dataf(!pipeline_dffe_13),
	.datag(gnd),
	.cin(\op_1~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~73_sumout ),
	.cout(\op_1~74 ),
	.shareout());
defparam \op_1~73 .extended_lut = "off";
defparam \op_1~73 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~73 .shared_arith = "off";

cyclonev_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_14),
	.datae(gnd),
	.dataf(!pipeline_dffe_14),
	.datag(gnd),
	.cin(\op_1~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

cyclonev_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_15),
	.datae(gnd),
	.dataf(!pipeline_dffe_15),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_16),
	.datae(gnd),
	.dataf(!pipeline_dffe_16),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_17),
	.datae(gnd),
	.dataf(!pipeline_dffe_17),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_18),
	.datae(gnd),
	.dataf(!pipeline_dffe_18),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_19),
	.datae(gnd),
	.dataf(!pipeline_dffe_19),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_20),
	.datae(gnd),
	.dataf(!pipeline_dffe_20),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_21),
	.datae(gnd),
	.dataf(!pipeline_dffe_21),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_22),
	.datae(gnd),
	.dataf(!pipeline_dffe_22),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_23),
	.datae(gnd),
	.dataf(!pipeline_dffe_23),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_24),
	.datae(gnd),
	.dataf(!pipeline_dffe_24),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_25),
	.datae(gnd),
	.dataf(!pipeline_dffe_25),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_26),
	.datae(gnd),
	.dataf(!pipeline_dffe_26),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_27),
	.datae(gnd),
	.dataf(!pipeline_dffe_27),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_28),
	.datae(gnd),
	.dataf(!pipeline_dffe_28),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

cyclonev_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_29),
	.datae(gnd),
	.dataf(!pipeline_dffe_29),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

cyclonev_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_30),
	.datae(gnd),
	.dataf(!pipeline_dffe_30),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

cyclonev_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_31),
	.datae(gnd),
	.dataf(!pipeline_dffe_31),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

endmodule

module sine_asj_dxx (
	dxxpdo_5,
	dxxpdo_6,
	dxxpdo_7,
	dxxpdo_8,
	dxxpdo_9,
	dxxpdo_10,
	dxxpdo_11,
	dxxpdo_12,
	dxxpdo_13,
	dxxpdo_14,
	dxxpdo_15,
	dxxpdo_16,
	dxxpdo_17,
	dxxpdo_20,
	dxxpdo_18,
	dxxpdo_19,
	dxxrv_3,
	dxxrv_2,
	dxxrv_1,
	dxxrv_0,
	data_out_12,
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_31,
	pipeline_dffe_15,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	NJQG9082,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dxxpdo_5;
output 	dxxpdo_6;
output 	dxxpdo_7;
output 	dxxpdo_8;
output 	dxxpdo_9;
output 	dxxpdo_10;
output 	dxxpdo_11;
output 	dxxpdo_12;
output 	dxxpdo_13;
output 	dxxpdo_14;
output 	dxxpdo_15;
output 	dxxpdo_16;
output 	dxxpdo_17;
output 	dxxpdo_20;
output 	dxxpdo_18;
output 	dxxpdo_19;
input 	dxxrv_3;
input 	dxxrv_2;
input 	dxxrv_1;
input 	dxxrv_0;
input 	data_out_12;
input 	pipeline_dffe_16;
input 	pipeline_dffe_17;
input 	pipeline_dffe_18;
input 	pipeline_dffe_19;
input 	pipeline_dffe_20;
input 	pipeline_dffe_21;
input 	pipeline_dffe_22;
input 	pipeline_dffe_23;
input 	pipeline_dffe_24;
input 	pipeline_dffe_25;
input 	pipeline_dffe_26;
input 	pipeline_dffe_27;
input 	pipeline_dffe_28;
input 	pipeline_dffe_31;
input 	pipeline_dffe_15;
input 	pipeline_dffe_29;
input 	pipeline_dffe_30;
input 	pipeline_dffe_14;
input 	pipeline_dffe_13;
input 	pipeline_dffe_12;
input 	pipeline_dffe_11;
input 	NJQG9082;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~82_cout ;
wire \Add0~78_cout ;
wire \Add0~74_cout ;
wire \Add0~70_cout ;
wire \Add0~58_cout ;
wire \Add0~1_sumout ;
wire \phi_dither_out_w[5]~q ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \phi_dither_out_w[6]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \phi_dither_out_w[7]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \phi_dither_out_w[8]~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \phi_dither_out_w[9]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \phi_dither_out_w[10]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \phi_dither_out_w[11]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \phi_dither_out_w[12]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \phi_dither_out_w[13]~q ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \phi_dither_out_w[14]~q ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \phi_dither_out_w[15]~q ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \phi_dither_out_w[16]~q ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \phi_dither_out_w[17]~q ;
wire \Add0~50 ;
wire \Add0~62 ;
wire \Add0~66 ;
wire \Add0~53_sumout ;
wire \phi_dither_out_w[20]~q ;
wire \Add0~61_sumout ;
wire \phi_dither_out_w[18]~q ;
wire \Add0~65_sumout ;
wire \phi_dither_out_w[19]~q ;


dffeas \dxxpdo[5] (
	.clk(clk),
	.d(\phi_dither_out_w[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_5),
	.prn(vcc));
defparam \dxxpdo[5] .is_wysiwyg = "true";
defparam \dxxpdo[5] .power_up = "low";

dffeas \dxxpdo[6] (
	.clk(clk),
	.d(\phi_dither_out_w[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_6),
	.prn(vcc));
defparam \dxxpdo[6] .is_wysiwyg = "true";
defparam \dxxpdo[6] .power_up = "low";

dffeas \dxxpdo[7] (
	.clk(clk),
	.d(\phi_dither_out_w[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_7),
	.prn(vcc));
defparam \dxxpdo[7] .is_wysiwyg = "true";
defparam \dxxpdo[7] .power_up = "low";

dffeas \dxxpdo[8] (
	.clk(clk),
	.d(\phi_dither_out_w[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_8),
	.prn(vcc));
defparam \dxxpdo[8] .is_wysiwyg = "true";
defparam \dxxpdo[8] .power_up = "low";

dffeas \dxxpdo[9] (
	.clk(clk),
	.d(\phi_dither_out_w[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_9),
	.prn(vcc));
defparam \dxxpdo[9] .is_wysiwyg = "true";
defparam \dxxpdo[9] .power_up = "low";

dffeas \dxxpdo[10] (
	.clk(clk),
	.d(\phi_dither_out_w[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_10),
	.prn(vcc));
defparam \dxxpdo[10] .is_wysiwyg = "true";
defparam \dxxpdo[10] .power_up = "low";

dffeas \dxxpdo[11] (
	.clk(clk),
	.d(\phi_dither_out_w[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_11),
	.prn(vcc));
defparam \dxxpdo[11] .is_wysiwyg = "true";
defparam \dxxpdo[11] .power_up = "low";

dffeas \dxxpdo[12] (
	.clk(clk),
	.d(\phi_dither_out_w[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_12),
	.prn(vcc));
defparam \dxxpdo[12] .is_wysiwyg = "true";
defparam \dxxpdo[12] .power_up = "low";

dffeas \dxxpdo[13] (
	.clk(clk),
	.d(\phi_dither_out_w[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_13),
	.prn(vcc));
defparam \dxxpdo[13] .is_wysiwyg = "true";
defparam \dxxpdo[13] .power_up = "low";

dffeas \dxxpdo[14] (
	.clk(clk),
	.d(\phi_dither_out_w[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_14),
	.prn(vcc));
defparam \dxxpdo[14] .is_wysiwyg = "true";
defparam \dxxpdo[14] .power_up = "low";

dffeas \dxxpdo[15] (
	.clk(clk),
	.d(\phi_dither_out_w[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_15),
	.prn(vcc));
defparam \dxxpdo[15] .is_wysiwyg = "true";
defparam \dxxpdo[15] .power_up = "low";

dffeas \dxxpdo[16] (
	.clk(clk),
	.d(\phi_dither_out_w[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_16),
	.prn(vcc));
defparam \dxxpdo[16] .is_wysiwyg = "true";
defparam \dxxpdo[16] .power_up = "low";

dffeas \dxxpdo[17] (
	.clk(clk),
	.d(\phi_dither_out_w[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_17),
	.prn(vcc));
defparam \dxxpdo[17] .is_wysiwyg = "true";
defparam \dxxpdo[17] .power_up = "low";

dffeas \dxxpdo[20] (
	.clk(clk),
	.d(\phi_dither_out_w[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_20),
	.prn(vcc));
defparam \dxxpdo[20] .is_wysiwyg = "true";
defparam \dxxpdo[20] .power_up = "low";

dffeas \dxxpdo[18] (
	.clk(clk),
	.d(\phi_dither_out_w[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_18),
	.prn(vcc));
defparam \dxxpdo[18] .is_wysiwyg = "true";
defparam \dxxpdo[18] .power_up = "low";

dffeas \dxxpdo[19] (
	.clk(clk),
	.d(\phi_dither_out_w[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxpdo_19),
	.prn(vcc));
defparam \dxxpdo[19] .is_wysiwyg = "true";
defparam \dxxpdo[19] .power_up = "low";

cyclonev_lcell_comb \Add0~82 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_0),
	.datae(gnd),
	.dataf(!pipeline_dffe_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~82_cout ),
	.shareout());
defparam \Add0~82 .extended_lut = "off";
defparam \Add0~82 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~82 .shared_arith = "off";

cyclonev_lcell_comb \Add0~78 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_1),
	.datae(gnd),
	.dataf(!pipeline_dffe_12),
	.datag(gnd),
	.cin(\Add0~82_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~78_cout ),
	.shareout());
defparam \Add0~78 .extended_lut = "off";
defparam \Add0~78 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~78 .shared_arith = "off";

cyclonev_lcell_comb \Add0~74 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_2),
	.datae(gnd),
	.dataf(!pipeline_dffe_13),
	.datag(gnd),
	.cin(\Add0~78_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~74_cout ),
	.shareout());
defparam \Add0~74 .extended_lut = "off";
defparam \Add0~74 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~74 .shared_arith = "off";

cyclonev_lcell_comb \Add0~70 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_14),
	.datag(gnd),
	.cin(\Add0~74_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~70_cout ),
	.shareout());
defparam \Add0~70 .extended_lut = "off";
defparam \Add0~70 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~70 .shared_arith = "off";

cyclonev_lcell_comb \Add0~58 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_15),
	.datag(gnd),
	.cin(\Add0~70_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~58_cout ),
	.shareout());
defparam \Add0~58 .extended_lut = "off";
defparam \Add0~58 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~58 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_16),
	.datag(gnd),
	.cin(\Add0~58_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \phi_dither_out_w[5] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[5]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[5] .is_wysiwyg = "true";
defparam \phi_dither_out_w[5] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_17),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \phi_dither_out_w[6] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[6]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[6] .is_wysiwyg = "true";
defparam \phi_dither_out_w[6] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_18),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \phi_dither_out_w[7] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[7]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[7] .is_wysiwyg = "true";
defparam \phi_dither_out_w[7] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_19),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \phi_dither_out_w[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[8]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[8] .is_wysiwyg = "true";
defparam \phi_dither_out_w[8] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_20),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \phi_dither_out_w[9] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[9]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[9] .is_wysiwyg = "true";
defparam \phi_dither_out_w[9] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_21),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \phi_dither_out_w[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[10]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[10] .is_wysiwyg = "true";
defparam \phi_dither_out_w[10] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_22),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \phi_dither_out_w[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[11]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[11] .is_wysiwyg = "true";
defparam \phi_dither_out_w[11] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_23),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \phi_dither_out_w[12] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[12]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[12] .is_wysiwyg = "true";
defparam \phi_dither_out_w[12] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_24),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \phi_dither_out_w[13] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[13]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[13] .is_wysiwyg = "true";
defparam \phi_dither_out_w[13] .power_up = "low";

cyclonev_lcell_comb \Add0~37 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_25),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \phi_dither_out_w[14] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[14]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[14] .is_wysiwyg = "true";
defparam \phi_dither_out_w[14] .power_up = "low";

cyclonev_lcell_comb \Add0~41 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_26),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \phi_dither_out_w[15] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[15]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[15] .is_wysiwyg = "true";
defparam \phi_dither_out_w[15] .power_up = "low";

cyclonev_lcell_comb \Add0~45 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_27),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \phi_dither_out_w[16] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[16]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[16] .is_wysiwyg = "true";
defparam \phi_dither_out_w[16] .power_up = "low";

cyclonev_lcell_comb \Add0~49 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_28),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~49 .shared_arith = "off";

dffeas \phi_dither_out_w[17] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[17]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[17] .is_wysiwyg = "true";
defparam \phi_dither_out_w[17] .power_up = "low";

cyclonev_lcell_comb \Add0~61 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_29),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~61 .shared_arith = "off";

cyclonev_lcell_comb \Add0~65 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_30),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~65 .shared_arith = "off";

cyclonev_lcell_comb \Add0~53 (
	.dataa(!NJQG9082),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_31),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF55000000FF;
defparam \Add0~53 .shared_arith = "off";

dffeas \phi_dither_out_w[20] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[20]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[20] .is_wysiwyg = "true";
defparam \phi_dither_out_w[20] .power_up = "low";

dffeas \phi_dither_out_w[18] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[18]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[18] .is_wysiwyg = "true";
defparam \phi_dither_out_w[18] .power_up = "low";

dffeas \phi_dither_out_w[19] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_dither_out_w[19]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[19] .is_wysiwyg = "true";
defparam \phi_dither_out_w[19] .power_up = "low";

endmodule

module sine_asj_dxx_g (
	dxxrv_3,
	dxxrv_2,
	dxxrv_1,
	dxxrv_0,
	data_out_12,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dxxrv_3;
output 	dxxrv_2;
output 	dxxrv_1;
output 	dxxrv_0;
input 	data_out_12;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lsfr_reg~10_combout ;
wire \lsfr_reg[0]~q ;
wire \lsfr_reg[1]~q ;
wire \lsfr_reg~9_combout ;
wire \lsfr_reg[2]~q ;
wire \lsfr_reg~8_combout ;
wire \lsfr_reg[3]~q ;
wire \lsfr_reg~7_combout ;
wire \lsfr_reg[4]~q ;
wire \lsfr_reg[5]~q ;
wire \lsfr_reg~6_combout ;
wire \lsfr_reg[6]~q ;
wire \lsfr_reg~5_combout ;
wire \lsfr_reg[7]~q ;
wire \lsfr_reg[8]~q ;
wire \lsfr_reg~3_combout ;
wire \lsfr_reg[9]~q ;
wire \lsfr_reg[10]~q ;
wire \lsfr_reg~2_combout ;
wire \lsfr_reg[11]~q ;
wire \lsfr_reg~1_combout ;
wire \lsfr_reg[12]~q ;
wire \lsfr_reg[13]~q ;
wire \lsfr_reg[14]~q ;
wire \lsfr_reg~0_combout ;
wire \lsfr_reg[15]~q ;
wire \Add0~0_combout ;
wire \Add0~1_combout ;
wire \Add0~2_combout ;
wire \lsfr_reg~4_combout ;


dffeas \dxxrv[3] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_3),
	.prn(vcc));
defparam \dxxrv[3] .is_wysiwyg = "true";
defparam \dxxrv[3] .power_up = "low";

dffeas \dxxrv[2] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_2),
	.prn(vcc));
defparam \dxxrv[2] .is_wysiwyg = "true";
defparam \dxxrv[2] .power_up = "low";

dffeas \dxxrv[1] (
	.clk(clk),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_1),
	.prn(vcc));
defparam \dxxrv[1] .is_wysiwyg = "true";
defparam \dxxrv[1] .power_up = "low";

dffeas \dxxrv[0] (
	.clk(clk),
	.d(\lsfr_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(dxxrv_0),
	.prn(vcc));
defparam \dxxrv[0] .is_wysiwyg = "true";
defparam \dxxrv[0] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~10 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[14]~q ),
	.datac(!\lsfr_reg[12]~q ),
	.datad(!\lsfr_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~10 .extended_lut = "off";
defparam \lsfr_reg~10 .lut_mask = 64'h6996699669966996;
defparam \lsfr_reg~10 .shared_arith = "off";

dffeas \lsfr_reg[0] (
	.clk(clk),
	.d(\lsfr_reg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(data_out_12),
	.q(\lsfr_reg[0]~q ),
	.prn(vcc));
defparam \lsfr_reg[0] .is_wysiwyg = "true";
defparam \lsfr_reg[0] .power_up = "low";

dffeas \lsfr_reg[1] (
	.clk(clk),
	.d(\lsfr_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[1]~q ),
	.prn(vcc));
defparam \lsfr_reg[1] .is_wysiwyg = "true";
defparam \lsfr_reg[1] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~9 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~9 .extended_lut = "off";
defparam \lsfr_reg~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~9 .shared_arith = "off";

dffeas \lsfr_reg[2] (
	.clk(clk),
	.d(\lsfr_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[2]~q ),
	.prn(vcc));
defparam \lsfr_reg[2] .is_wysiwyg = "true";
defparam \lsfr_reg[2] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~8 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~8 .extended_lut = "off";
defparam \lsfr_reg~8 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~8 .shared_arith = "off";

dffeas \lsfr_reg[3] (
	.clk(clk),
	.d(\lsfr_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[3]~q ),
	.prn(vcc));
defparam \lsfr_reg[3] .is_wysiwyg = "true";
defparam \lsfr_reg[3] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~7 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~7 .extended_lut = "off";
defparam \lsfr_reg~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~7 .shared_arith = "off";

dffeas \lsfr_reg[4] (
	.clk(clk),
	.d(\lsfr_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[4]~q ),
	.prn(vcc));
defparam \lsfr_reg[4] .is_wysiwyg = "true";
defparam \lsfr_reg[4] .power_up = "low";

dffeas \lsfr_reg[5] (
	.clk(clk),
	.d(\lsfr_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[5]~q ),
	.prn(vcc));
defparam \lsfr_reg[5] .is_wysiwyg = "true";
defparam \lsfr_reg[5] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~6 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~6 .extended_lut = "off";
defparam \lsfr_reg~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~6 .shared_arith = "off";

dffeas \lsfr_reg[6] (
	.clk(clk),
	.d(\lsfr_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[6]~q ),
	.prn(vcc));
defparam \lsfr_reg[6] .is_wysiwyg = "true";
defparam \lsfr_reg[6] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~5 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~5 .extended_lut = "off";
defparam \lsfr_reg~5 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~5 .shared_arith = "off";

dffeas \lsfr_reg[7] (
	.clk(clk),
	.d(\lsfr_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[7]~q ),
	.prn(vcc));
defparam \lsfr_reg[7] .is_wysiwyg = "true";
defparam \lsfr_reg[7] .power_up = "low";

dffeas \lsfr_reg[8] (
	.clk(clk),
	.d(\lsfr_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[8]~q ),
	.prn(vcc));
defparam \lsfr_reg[8] .is_wysiwyg = "true";
defparam \lsfr_reg[8] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~3 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~3 .extended_lut = "off";
defparam \lsfr_reg~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~3 .shared_arith = "off";

dffeas \lsfr_reg[9] (
	.clk(clk),
	.d(\lsfr_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[9]~q ),
	.prn(vcc));
defparam \lsfr_reg[9] .is_wysiwyg = "true";
defparam \lsfr_reg[9] .power_up = "low";

dffeas \lsfr_reg[10] (
	.clk(clk),
	.d(\lsfr_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[10]~q ),
	.prn(vcc));
defparam \lsfr_reg[10] .is_wysiwyg = "true";
defparam \lsfr_reg[10] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~2 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~2 .extended_lut = "off";
defparam \lsfr_reg~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~2 .shared_arith = "off";

dffeas \lsfr_reg[11] (
	.clk(clk),
	.d(\lsfr_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[11]~q ),
	.prn(vcc));
defparam \lsfr_reg[11] .is_wysiwyg = "true";
defparam \lsfr_reg[11] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~1 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~1 .extended_lut = "off";
defparam \lsfr_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~1 .shared_arith = "off";

dffeas \lsfr_reg[12] (
	.clk(clk),
	.d(\lsfr_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[12]~q ),
	.prn(vcc));
defparam \lsfr_reg[12] .is_wysiwyg = "true";
defparam \lsfr_reg[12] .power_up = "low";

dffeas \lsfr_reg[13] (
	.clk(clk),
	.d(\lsfr_reg[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[13]~q ),
	.prn(vcc));
defparam \lsfr_reg[13] .is_wysiwyg = "true";
defparam \lsfr_reg[13] .power_up = "low";

dffeas \lsfr_reg[14] (
	.clk(clk),
	.d(\lsfr_reg[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[14]~q ),
	.prn(vcc));
defparam \lsfr_reg[14] .is_wysiwyg = "true";
defparam \lsfr_reg[14] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~0 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~0 .extended_lut = "off";
defparam \lsfr_reg~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~0 .shared_arith = "off";

dffeas \lsfr_reg[15] (
	.clk(clk),
	.d(\lsfr_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_out_12),
	.q(\lsfr_reg[15]~q ),
	.prn(vcc));
defparam \lsfr_reg[15] .is_wysiwyg = "true";
defparam \lsfr_reg[15] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[14]~q ),
	.datac(!\lsfr_reg[13]~q ),
	.datad(!\lsfr_reg[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[14]~q ),
	.datac(!\lsfr_reg[13]~q ),
	.datad(!\lsfr_reg[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6996699669966996;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[13]~q ),
	.datac(!\lsfr_reg[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h9696969696969696;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \lsfr_reg~4 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~4 .extended_lut = "off";
defparam \lsfr_reg~4 .lut_mask = 64'h6666666666666666;
defparam \lsfr_reg~4 .shared_arith = "off";

endmodule

module sine_asj_gal (
	rom_add_0,
	rom_add_1,
	rom_add_2,
	rom_add_3,
	rom_add_4,
	rom_add_5,
	rom_add_6,
	rom_add_7,
	rom_add_8,
	rom_add_9,
	rom_add_10,
	rom_add_11,
	rom_add_12,
	rom_add_15,
	rom_add_13,
	rom_add_14,
	data_out_12,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_15,
	pipeline_dffe_13,
	pipeline_dffe_14,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	rom_add_0;
output 	rom_add_1;
output 	rom_add_2;
output 	rom_add_3;
output 	rom_add_4;
output 	rom_add_5;
output 	rom_add_6;
output 	rom_add_7;
output 	rom_add_8;
output 	rom_add_9;
output 	rom_add_10;
output 	rom_add_11;
output 	rom_add_12;
output 	rom_add_15;
output 	rom_add_13;
output 	rom_add_14;
input 	data_out_12;
input 	pipeline_dffe_0;
input 	pipeline_dffe_1;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	pipeline_dffe_12;
input 	pipeline_dffe_15;
input 	pipeline_dffe_13;
input 	pipeline_dffe_14;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \rom_add[0] (
	.clk(clk),
	.d(pipeline_dffe_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_0),
	.prn(vcc));
defparam \rom_add[0] .is_wysiwyg = "true";
defparam \rom_add[0] .power_up = "low";

dffeas \rom_add[1] (
	.clk(clk),
	.d(pipeline_dffe_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_1),
	.prn(vcc));
defparam \rom_add[1] .is_wysiwyg = "true";
defparam \rom_add[1] .power_up = "low";

dffeas \rom_add[2] (
	.clk(clk),
	.d(pipeline_dffe_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_2),
	.prn(vcc));
defparam \rom_add[2] .is_wysiwyg = "true";
defparam \rom_add[2] .power_up = "low";

dffeas \rom_add[3] (
	.clk(clk),
	.d(pipeline_dffe_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_3),
	.prn(vcc));
defparam \rom_add[3] .is_wysiwyg = "true";
defparam \rom_add[3] .power_up = "low";

dffeas \rom_add[4] (
	.clk(clk),
	.d(pipeline_dffe_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_4),
	.prn(vcc));
defparam \rom_add[4] .is_wysiwyg = "true";
defparam \rom_add[4] .power_up = "low";

dffeas \rom_add[5] (
	.clk(clk),
	.d(pipeline_dffe_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_5),
	.prn(vcc));
defparam \rom_add[5] .is_wysiwyg = "true";
defparam \rom_add[5] .power_up = "low";

dffeas \rom_add[6] (
	.clk(clk),
	.d(pipeline_dffe_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_6),
	.prn(vcc));
defparam \rom_add[6] .is_wysiwyg = "true";
defparam \rom_add[6] .power_up = "low";

dffeas \rom_add[7] (
	.clk(clk),
	.d(pipeline_dffe_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_7),
	.prn(vcc));
defparam \rom_add[7] .is_wysiwyg = "true";
defparam \rom_add[7] .power_up = "low";

dffeas \rom_add[8] (
	.clk(clk),
	.d(pipeline_dffe_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_8),
	.prn(vcc));
defparam \rom_add[8] .is_wysiwyg = "true";
defparam \rom_add[8] .power_up = "low";

dffeas \rom_add[9] (
	.clk(clk),
	.d(pipeline_dffe_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_9),
	.prn(vcc));
defparam \rom_add[9] .is_wysiwyg = "true";
defparam \rom_add[9] .power_up = "low";

dffeas \rom_add[10] (
	.clk(clk),
	.d(pipeline_dffe_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_10),
	.prn(vcc));
defparam \rom_add[10] .is_wysiwyg = "true";
defparam \rom_add[10] .power_up = "low";

dffeas \rom_add[11] (
	.clk(clk),
	.d(pipeline_dffe_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_11),
	.prn(vcc));
defparam \rom_add[11] .is_wysiwyg = "true";
defparam \rom_add[11] .power_up = "low";

dffeas \rom_add[12] (
	.clk(clk),
	.d(pipeline_dffe_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_12),
	.prn(vcc));
defparam \rom_add[12] .is_wysiwyg = "true";
defparam \rom_add[12] .power_up = "low";

dffeas \rom_add[15] (
	.clk(clk),
	.d(pipeline_dffe_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_15),
	.prn(vcc));
defparam \rom_add[15] .is_wysiwyg = "true";
defparam \rom_add[15] .power_up = "low";

dffeas \rom_add[13] (
	.clk(clk),
	.d(pipeline_dffe_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_13),
	.prn(vcc));
defparam \rom_add[13] .is_wysiwyg = "true";
defparam \rom_add[13] .power_up = "low";

dffeas \rom_add[14] (
	.clk(clk),
	.d(pipeline_dffe_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(rom_add_14),
	.prn(vcc));
defparam \rom_add[14] .is_wysiwyg = "true";
defparam \rom_add[14] .power_up = "low";

endmodule

module sine_asj_nco_as_m_cen (
	ram_block1a96,
	ram_block1a120,
	ram_block1a144,
	ram_block1a168,
	ram_block1a48,
	ram_block1a72,
	ram_block1a0,
	ram_block1a24,
	ram_block1a97,
	ram_block1a121,
	ram_block1a145,
	ram_block1a169,
	ram_block1a49,
	ram_block1a73,
	ram_block1a1,
	ram_block1a25,
	ram_block1a98,
	ram_block1a122,
	ram_block1a146,
	ram_block1a170,
	ram_block1a50,
	ram_block1a74,
	ram_block1a2,
	ram_block1a26,
	ram_block1a99,
	ram_block1a123,
	ram_block1a147,
	ram_block1a171,
	ram_block1a51,
	ram_block1a75,
	ram_block1a3,
	ram_block1a27,
	ram_block1a100,
	ram_block1a124,
	ram_block1a148,
	ram_block1a172,
	ram_block1a52,
	ram_block1a76,
	ram_block1a4,
	ram_block1a28,
	ram_block1a101,
	ram_block1a125,
	ram_block1a149,
	ram_block1a173,
	ram_block1a53,
	ram_block1a77,
	ram_block1a5,
	ram_block1a29,
	ram_block1a102,
	ram_block1a126,
	ram_block1a150,
	ram_block1a174,
	ram_block1a54,
	ram_block1a78,
	ram_block1a6,
	ram_block1a30,
	ram_block1a103,
	ram_block1a127,
	ram_block1a151,
	ram_block1a175,
	ram_block1a55,
	ram_block1a79,
	ram_block1a7,
	ram_block1a31,
	ram_block1a104,
	ram_block1a128,
	ram_block1a152,
	ram_block1a176,
	ram_block1a56,
	ram_block1a80,
	ram_block1a8,
	ram_block1a32,
	ram_block1a105,
	ram_block1a129,
	ram_block1a153,
	ram_block1a177,
	ram_block1a57,
	ram_block1a81,
	ram_block1a9,
	ram_block1a33,
	ram_block1a106,
	ram_block1a130,
	ram_block1a154,
	ram_block1a178,
	ram_block1a58,
	ram_block1a82,
	ram_block1a10,
	ram_block1a34,
	ram_block1a107,
	ram_block1a131,
	ram_block1a155,
	ram_block1a179,
	ram_block1a59,
	ram_block1a83,
	ram_block1a11,
	ram_block1a35,
	ram_block1a108,
	ram_block1a132,
	ram_block1a156,
	ram_block1a180,
	ram_block1a60,
	ram_block1a84,
	ram_block1a12,
	ram_block1a36,
	ram_block1a109,
	ram_block1a133,
	ram_block1a157,
	ram_block1a181,
	ram_block1a61,
	ram_block1a85,
	ram_block1a13,
	ram_block1a37,
	ram_block1a110,
	ram_block1a134,
	ram_block1a158,
	ram_block1a182,
	ram_block1a62,
	ram_block1a86,
	ram_block1a14,
	ram_block1a38,
	ram_block1a111,
	ram_block1a135,
	ram_block1a159,
	ram_block1a183,
	ram_block1a63,
	ram_block1a87,
	ram_block1a15,
	ram_block1a39,
	ram_block1a112,
	ram_block1a136,
	ram_block1a160,
	ram_block1a184,
	ram_block1a64,
	ram_block1a88,
	ram_block1a16,
	ram_block1a40,
	ram_block1a113,
	ram_block1a137,
	ram_block1a161,
	ram_block1a185,
	ram_block1a65,
	ram_block1a89,
	ram_block1a17,
	ram_block1a41,
	ram_block1a114,
	ram_block1a138,
	ram_block1a162,
	ram_block1a186,
	ram_block1a66,
	ram_block1a90,
	ram_block1a18,
	ram_block1a42,
	ram_block1a115,
	ram_block1a139,
	ram_block1a163,
	ram_block1a187,
	ram_block1a67,
	ram_block1a91,
	ram_block1a19,
	ram_block1a43,
	ram_block1a116,
	ram_block1a140,
	ram_block1a164,
	ram_block1a188,
	ram_block1a68,
	ram_block1a92,
	ram_block1a20,
	ram_block1a44,
	ram_block1a117,
	ram_block1a141,
	ram_block1a165,
	ram_block1a189,
	ram_block1a69,
	ram_block1a93,
	ram_block1a21,
	ram_block1a45,
	ram_block1a118,
	ram_block1a142,
	ram_block1a166,
	ram_block1a190,
	ram_block1a70,
	ram_block1a94,
	ram_block1a22,
	ram_block1a46,
	ram_block1a119,
	ram_block1a143,
	ram_block1a167,
	ram_block1a191,
	ram_block1a71,
	ram_block1a95,
	ram_block1a23,
	ram_block1a47,
	rom_add_0,
	rom_add_1,
	rom_add_2,
	rom_add_3,
	rom_add_4,
	rom_add_5,
	rom_add_6,
	rom_add_7,
	rom_add_8,
	rom_add_9,
	rom_add_10,
	rom_add_11,
	rom_add_12,
	rom_add_15,
	rom_add_13,
	rom_add_14,
	out_address_reg_a_2,
	out_address_reg_a_0,
	out_address_reg_a_1,
	clk,
	clken)/* synthesis synthesis_greybox=1 */;
output 	ram_block1a96;
output 	ram_block1a120;
output 	ram_block1a144;
output 	ram_block1a168;
output 	ram_block1a48;
output 	ram_block1a72;
output 	ram_block1a0;
output 	ram_block1a24;
output 	ram_block1a97;
output 	ram_block1a121;
output 	ram_block1a145;
output 	ram_block1a169;
output 	ram_block1a49;
output 	ram_block1a73;
output 	ram_block1a1;
output 	ram_block1a25;
output 	ram_block1a98;
output 	ram_block1a122;
output 	ram_block1a146;
output 	ram_block1a170;
output 	ram_block1a50;
output 	ram_block1a74;
output 	ram_block1a2;
output 	ram_block1a26;
output 	ram_block1a99;
output 	ram_block1a123;
output 	ram_block1a147;
output 	ram_block1a171;
output 	ram_block1a51;
output 	ram_block1a75;
output 	ram_block1a3;
output 	ram_block1a27;
output 	ram_block1a100;
output 	ram_block1a124;
output 	ram_block1a148;
output 	ram_block1a172;
output 	ram_block1a52;
output 	ram_block1a76;
output 	ram_block1a4;
output 	ram_block1a28;
output 	ram_block1a101;
output 	ram_block1a125;
output 	ram_block1a149;
output 	ram_block1a173;
output 	ram_block1a53;
output 	ram_block1a77;
output 	ram_block1a5;
output 	ram_block1a29;
output 	ram_block1a102;
output 	ram_block1a126;
output 	ram_block1a150;
output 	ram_block1a174;
output 	ram_block1a54;
output 	ram_block1a78;
output 	ram_block1a6;
output 	ram_block1a30;
output 	ram_block1a103;
output 	ram_block1a127;
output 	ram_block1a151;
output 	ram_block1a175;
output 	ram_block1a55;
output 	ram_block1a79;
output 	ram_block1a7;
output 	ram_block1a31;
output 	ram_block1a104;
output 	ram_block1a128;
output 	ram_block1a152;
output 	ram_block1a176;
output 	ram_block1a56;
output 	ram_block1a80;
output 	ram_block1a8;
output 	ram_block1a32;
output 	ram_block1a105;
output 	ram_block1a129;
output 	ram_block1a153;
output 	ram_block1a177;
output 	ram_block1a57;
output 	ram_block1a81;
output 	ram_block1a9;
output 	ram_block1a33;
output 	ram_block1a106;
output 	ram_block1a130;
output 	ram_block1a154;
output 	ram_block1a178;
output 	ram_block1a58;
output 	ram_block1a82;
output 	ram_block1a10;
output 	ram_block1a34;
output 	ram_block1a107;
output 	ram_block1a131;
output 	ram_block1a155;
output 	ram_block1a179;
output 	ram_block1a59;
output 	ram_block1a83;
output 	ram_block1a11;
output 	ram_block1a35;
output 	ram_block1a108;
output 	ram_block1a132;
output 	ram_block1a156;
output 	ram_block1a180;
output 	ram_block1a60;
output 	ram_block1a84;
output 	ram_block1a12;
output 	ram_block1a36;
output 	ram_block1a109;
output 	ram_block1a133;
output 	ram_block1a157;
output 	ram_block1a181;
output 	ram_block1a61;
output 	ram_block1a85;
output 	ram_block1a13;
output 	ram_block1a37;
output 	ram_block1a110;
output 	ram_block1a134;
output 	ram_block1a158;
output 	ram_block1a182;
output 	ram_block1a62;
output 	ram_block1a86;
output 	ram_block1a14;
output 	ram_block1a38;
output 	ram_block1a111;
output 	ram_block1a135;
output 	ram_block1a159;
output 	ram_block1a183;
output 	ram_block1a63;
output 	ram_block1a87;
output 	ram_block1a15;
output 	ram_block1a39;
output 	ram_block1a112;
output 	ram_block1a136;
output 	ram_block1a160;
output 	ram_block1a184;
output 	ram_block1a64;
output 	ram_block1a88;
output 	ram_block1a16;
output 	ram_block1a40;
output 	ram_block1a113;
output 	ram_block1a137;
output 	ram_block1a161;
output 	ram_block1a185;
output 	ram_block1a65;
output 	ram_block1a89;
output 	ram_block1a17;
output 	ram_block1a41;
output 	ram_block1a114;
output 	ram_block1a138;
output 	ram_block1a162;
output 	ram_block1a186;
output 	ram_block1a66;
output 	ram_block1a90;
output 	ram_block1a18;
output 	ram_block1a42;
output 	ram_block1a115;
output 	ram_block1a139;
output 	ram_block1a163;
output 	ram_block1a187;
output 	ram_block1a67;
output 	ram_block1a91;
output 	ram_block1a19;
output 	ram_block1a43;
output 	ram_block1a116;
output 	ram_block1a140;
output 	ram_block1a164;
output 	ram_block1a188;
output 	ram_block1a68;
output 	ram_block1a92;
output 	ram_block1a20;
output 	ram_block1a44;
output 	ram_block1a117;
output 	ram_block1a141;
output 	ram_block1a165;
output 	ram_block1a189;
output 	ram_block1a69;
output 	ram_block1a93;
output 	ram_block1a21;
output 	ram_block1a45;
output 	ram_block1a118;
output 	ram_block1a142;
output 	ram_block1a166;
output 	ram_block1a190;
output 	ram_block1a70;
output 	ram_block1a94;
output 	ram_block1a22;
output 	ram_block1a46;
output 	ram_block1a119;
output 	ram_block1a143;
output 	ram_block1a167;
output 	ram_block1a191;
output 	ram_block1a71;
output 	ram_block1a95;
output 	ram_block1a23;
output 	ram_block1a47;
input 	rom_add_0;
input 	rom_add_1;
input 	rom_add_2;
input 	rom_add_3;
input 	rom_add_4;
input 	rom_add_5;
input 	rom_add_6;
input 	rom_add_7;
input 	rom_add_8;
input 	rom_add_9;
input 	rom_add_10;
input 	rom_add_11;
input 	rom_add_12;
input 	rom_add_15;
input 	rom_add_13;
input 	rom_add_14;
output 	out_address_reg_a_2;
output 	out_address_reg_a_0;
output 	out_address_reg_a_1;
input 	clk;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_altsyncram_1 altsyncram_component0(
	.ram_block1a96(ram_block1a96),
	.ram_block1a120(ram_block1a120),
	.ram_block1a144(ram_block1a144),
	.ram_block1a168(ram_block1a168),
	.ram_block1a48(ram_block1a48),
	.ram_block1a72(ram_block1a72),
	.ram_block1a0(ram_block1a0),
	.ram_block1a24(ram_block1a24),
	.ram_block1a97(ram_block1a97),
	.ram_block1a121(ram_block1a121),
	.ram_block1a145(ram_block1a145),
	.ram_block1a169(ram_block1a169),
	.ram_block1a49(ram_block1a49),
	.ram_block1a73(ram_block1a73),
	.ram_block1a1(ram_block1a1),
	.ram_block1a25(ram_block1a25),
	.ram_block1a98(ram_block1a98),
	.ram_block1a122(ram_block1a122),
	.ram_block1a146(ram_block1a146),
	.ram_block1a170(ram_block1a170),
	.ram_block1a50(ram_block1a50),
	.ram_block1a74(ram_block1a74),
	.ram_block1a2(ram_block1a2),
	.ram_block1a26(ram_block1a26),
	.ram_block1a99(ram_block1a99),
	.ram_block1a123(ram_block1a123),
	.ram_block1a147(ram_block1a147),
	.ram_block1a171(ram_block1a171),
	.ram_block1a51(ram_block1a51),
	.ram_block1a75(ram_block1a75),
	.ram_block1a3(ram_block1a3),
	.ram_block1a27(ram_block1a27),
	.ram_block1a100(ram_block1a100),
	.ram_block1a124(ram_block1a124),
	.ram_block1a148(ram_block1a148),
	.ram_block1a172(ram_block1a172),
	.ram_block1a52(ram_block1a52),
	.ram_block1a76(ram_block1a76),
	.ram_block1a4(ram_block1a4),
	.ram_block1a28(ram_block1a28),
	.ram_block1a101(ram_block1a101),
	.ram_block1a125(ram_block1a125),
	.ram_block1a149(ram_block1a149),
	.ram_block1a173(ram_block1a173),
	.ram_block1a53(ram_block1a53),
	.ram_block1a77(ram_block1a77),
	.ram_block1a5(ram_block1a5),
	.ram_block1a29(ram_block1a29),
	.ram_block1a102(ram_block1a102),
	.ram_block1a126(ram_block1a126),
	.ram_block1a150(ram_block1a150),
	.ram_block1a174(ram_block1a174),
	.ram_block1a54(ram_block1a54),
	.ram_block1a78(ram_block1a78),
	.ram_block1a6(ram_block1a6),
	.ram_block1a30(ram_block1a30),
	.ram_block1a103(ram_block1a103),
	.ram_block1a127(ram_block1a127),
	.ram_block1a151(ram_block1a151),
	.ram_block1a175(ram_block1a175),
	.ram_block1a55(ram_block1a55),
	.ram_block1a79(ram_block1a79),
	.ram_block1a7(ram_block1a7),
	.ram_block1a31(ram_block1a31),
	.ram_block1a104(ram_block1a104),
	.ram_block1a128(ram_block1a128),
	.ram_block1a152(ram_block1a152),
	.ram_block1a176(ram_block1a176),
	.ram_block1a56(ram_block1a56),
	.ram_block1a80(ram_block1a80),
	.ram_block1a8(ram_block1a8),
	.ram_block1a32(ram_block1a32),
	.ram_block1a105(ram_block1a105),
	.ram_block1a129(ram_block1a129),
	.ram_block1a153(ram_block1a153),
	.ram_block1a177(ram_block1a177),
	.ram_block1a57(ram_block1a57),
	.ram_block1a81(ram_block1a81),
	.ram_block1a9(ram_block1a9),
	.ram_block1a33(ram_block1a33),
	.ram_block1a106(ram_block1a106),
	.ram_block1a130(ram_block1a130),
	.ram_block1a154(ram_block1a154),
	.ram_block1a178(ram_block1a178),
	.ram_block1a58(ram_block1a58),
	.ram_block1a82(ram_block1a82),
	.ram_block1a10(ram_block1a10),
	.ram_block1a34(ram_block1a34),
	.ram_block1a107(ram_block1a107),
	.ram_block1a131(ram_block1a131),
	.ram_block1a155(ram_block1a155),
	.ram_block1a179(ram_block1a179),
	.ram_block1a59(ram_block1a59),
	.ram_block1a83(ram_block1a83),
	.ram_block1a11(ram_block1a11),
	.ram_block1a35(ram_block1a35),
	.ram_block1a108(ram_block1a108),
	.ram_block1a132(ram_block1a132),
	.ram_block1a156(ram_block1a156),
	.ram_block1a180(ram_block1a180),
	.ram_block1a60(ram_block1a60),
	.ram_block1a84(ram_block1a84),
	.ram_block1a12(ram_block1a12),
	.ram_block1a36(ram_block1a36),
	.ram_block1a109(ram_block1a109),
	.ram_block1a133(ram_block1a133),
	.ram_block1a157(ram_block1a157),
	.ram_block1a181(ram_block1a181),
	.ram_block1a61(ram_block1a61),
	.ram_block1a85(ram_block1a85),
	.ram_block1a13(ram_block1a13),
	.ram_block1a37(ram_block1a37),
	.ram_block1a110(ram_block1a110),
	.ram_block1a134(ram_block1a134),
	.ram_block1a158(ram_block1a158),
	.ram_block1a182(ram_block1a182),
	.ram_block1a62(ram_block1a62),
	.ram_block1a86(ram_block1a86),
	.ram_block1a14(ram_block1a14),
	.ram_block1a38(ram_block1a38),
	.ram_block1a111(ram_block1a111),
	.ram_block1a135(ram_block1a135),
	.ram_block1a159(ram_block1a159),
	.ram_block1a183(ram_block1a183),
	.ram_block1a63(ram_block1a63),
	.ram_block1a87(ram_block1a87),
	.ram_block1a15(ram_block1a15),
	.ram_block1a39(ram_block1a39),
	.ram_block1a112(ram_block1a112),
	.ram_block1a136(ram_block1a136),
	.ram_block1a160(ram_block1a160),
	.ram_block1a184(ram_block1a184),
	.ram_block1a64(ram_block1a64),
	.ram_block1a88(ram_block1a88),
	.ram_block1a16(ram_block1a16),
	.ram_block1a40(ram_block1a40),
	.ram_block1a113(ram_block1a113),
	.ram_block1a137(ram_block1a137),
	.ram_block1a161(ram_block1a161),
	.ram_block1a185(ram_block1a185),
	.ram_block1a65(ram_block1a65),
	.ram_block1a89(ram_block1a89),
	.ram_block1a17(ram_block1a17),
	.ram_block1a41(ram_block1a41),
	.ram_block1a114(ram_block1a114),
	.ram_block1a138(ram_block1a138),
	.ram_block1a162(ram_block1a162),
	.ram_block1a186(ram_block1a186),
	.ram_block1a66(ram_block1a66),
	.ram_block1a90(ram_block1a90),
	.ram_block1a18(ram_block1a18),
	.ram_block1a42(ram_block1a42),
	.ram_block1a115(ram_block1a115),
	.ram_block1a139(ram_block1a139),
	.ram_block1a163(ram_block1a163),
	.ram_block1a187(ram_block1a187),
	.ram_block1a67(ram_block1a67),
	.ram_block1a91(ram_block1a91),
	.ram_block1a19(ram_block1a19),
	.ram_block1a43(ram_block1a43),
	.ram_block1a116(ram_block1a116),
	.ram_block1a140(ram_block1a140),
	.ram_block1a164(ram_block1a164),
	.ram_block1a188(ram_block1a188),
	.ram_block1a68(ram_block1a68),
	.ram_block1a92(ram_block1a92),
	.ram_block1a20(ram_block1a20),
	.ram_block1a44(ram_block1a44),
	.ram_block1a117(ram_block1a117),
	.ram_block1a141(ram_block1a141),
	.ram_block1a165(ram_block1a165),
	.ram_block1a189(ram_block1a189),
	.ram_block1a69(ram_block1a69),
	.ram_block1a93(ram_block1a93),
	.ram_block1a21(ram_block1a21),
	.ram_block1a45(ram_block1a45),
	.ram_block1a118(ram_block1a118),
	.ram_block1a142(ram_block1a142),
	.ram_block1a166(ram_block1a166),
	.ram_block1a190(ram_block1a190),
	.ram_block1a70(ram_block1a70),
	.ram_block1a94(ram_block1a94),
	.ram_block1a22(ram_block1a22),
	.ram_block1a46(ram_block1a46),
	.ram_block1a119(ram_block1a119),
	.ram_block1a143(ram_block1a143),
	.ram_block1a167(ram_block1a167),
	.ram_block1a191(ram_block1a191),
	.ram_block1a71(ram_block1a71),
	.ram_block1a95(ram_block1a95),
	.ram_block1a23(ram_block1a23),
	.ram_block1a47(ram_block1a47),
	.address_a({rom_add_15,rom_add_14,rom_add_13,rom_add_12,rom_add_11,rom_add_10,rom_add_9,rom_add_8,rom_add_7,rom_add_6,rom_add_5,rom_add_4,rom_add_3,rom_add_2,rom_add_1,rom_add_0}),
	.out_address_reg_a_2(out_address_reg_a_2),
	.out_address_reg_a_0(out_address_reg_a_0),
	.out_address_reg_a_1(out_address_reg_a_1),
	.clock0(clk),
	.clocken0(clken));

endmodule

module sine_altsyncram_1 (
	ram_block1a96,
	ram_block1a120,
	ram_block1a144,
	ram_block1a168,
	ram_block1a48,
	ram_block1a72,
	ram_block1a0,
	ram_block1a24,
	ram_block1a97,
	ram_block1a121,
	ram_block1a145,
	ram_block1a169,
	ram_block1a49,
	ram_block1a73,
	ram_block1a1,
	ram_block1a25,
	ram_block1a98,
	ram_block1a122,
	ram_block1a146,
	ram_block1a170,
	ram_block1a50,
	ram_block1a74,
	ram_block1a2,
	ram_block1a26,
	ram_block1a99,
	ram_block1a123,
	ram_block1a147,
	ram_block1a171,
	ram_block1a51,
	ram_block1a75,
	ram_block1a3,
	ram_block1a27,
	ram_block1a100,
	ram_block1a124,
	ram_block1a148,
	ram_block1a172,
	ram_block1a52,
	ram_block1a76,
	ram_block1a4,
	ram_block1a28,
	ram_block1a101,
	ram_block1a125,
	ram_block1a149,
	ram_block1a173,
	ram_block1a53,
	ram_block1a77,
	ram_block1a5,
	ram_block1a29,
	ram_block1a102,
	ram_block1a126,
	ram_block1a150,
	ram_block1a174,
	ram_block1a54,
	ram_block1a78,
	ram_block1a6,
	ram_block1a30,
	ram_block1a103,
	ram_block1a127,
	ram_block1a151,
	ram_block1a175,
	ram_block1a55,
	ram_block1a79,
	ram_block1a7,
	ram_block1a31,
	ram_block1a104,
	ram_block1a128,
	ram_block1a152,
	ram_block1a176,
	ram_block1a56,
	ram_block1a80,
	ram_block1a8,
	ram_block1a32,
	ram_block1a105,
	ram_block1a129,
	ram_block1a153,
	ram_block1a177,
	ram_block1a57,
	ram_block1a81,
	ram_block1a9,
	ram_block1a33,
	ram_block1a106,
	ram_block1a130,
	ram_block1a154,
	ram_block1a178,
	ram_block1a58,
	ram_block1a82,
	ram_block1a10,
	ram_block1a34,
	ram_block1a107,
	ram_block1a131,
	ram_block1a155,
	ram_block1a179,
	ram_block1a59,
	ram_block1a83,
	ram_block1a11,
	ram_block1a35,
	ram_block1a108,
	ram_block1a132,
	ram_block1a156,
	ram_block1a180,
	ram_block1a60,
	ram_block1a84,
	ram_block1a12,
	ram_block1a36,
	ram_block1a109,
	ram_block1a133,
	ram_block1a157,
	ram_block1a181,
	ram_block1a61,
	ram_block1a85,
	ram_block1a13,
	ram_block1a37,
	ram_block1a110,
	ram_block1a134,
	ram_block1a158,
	ram_block1a182,
	ram_block1a62,
	ram_block1a86,
	ram_block1a14,
	ram_block1a38,
	ram_block1a111,
	ram_block1a135,
	ram_block1a159,
	ram_block1a183,
	ram_block1a63,
	ram_block1a87,
	ram_block1a15,
	ram_block1a39,
	ram_block1a112,
	ram_block1a136,
	ram_block1a160,
	ram_block1a184,
	ram_block1a64,
	ram_block1a88,
	ram_block1a16,
	ram_block1a40,
	ram_block1a113,
	ram_block1a137,
	ram_block1a161,
	ram_block1a185,
	ram_block1a65,
	ram_block1a89,
	ram_block1a17,
	ram_block1a41,
	ram_block1a114,
	ram_block1a138,
	ram_block1a162,
	ram_block1a186,
	ram_block1a66,
	ram_block1a90,
	ram_block1a18,
	ram_block1a42,
	ram_block1a115,
	ram_block1a139,
	ram_block1a163,
	ram_block1a187,
	ram_block1a67,
	ram_block1a91,
	ram_block1a19,
	ram_block1a43,
	ram_block1a116,
	ram_block1a140,
	ram_block1a164,
	ram_block1a188,
	ram_block1a68,
	ram_block1a92,
	ram_block1a20,
	ram_block1a44,
	ram_block1a117,
	ram_block1a141,
	ram_block1a165,
	ram_block1a189,
	ram_block1a69,
	ram_block1a93,
	ram_block1a21,
	ram_block1a45,
	ram_block1a118,
	ram_block1a142,
	ram_block1a166,
	ram_block1a190,
	ram_block1a70,
	ram_block1a94,
	ram_block1a22,
	ram_block1a46,
	ram_block1a119,
	ram_block1a143,
	ram_block1a167,
	ram_block1a191,
	ram_block1a71,
	ram_block1a95,
	ram_block1a23,
	ram_block1a47,
	address_a,
	out_address_reg_a_2,
	out_address_reg_a_0,
	out_address_reg_a_1,
	clock0,
	clocken0)/* synthesis synthesis_greybox=1 */;
output 	ram_block1a96;
output 	ram_block1a120;
output 	ram_block1a144;
output 	ram_block1a168;
output 	ram_block1a48;
output 	ram_block1a72;
output 	ram_block1a0;
output 	ram_block1a24;
output 	ram_block1a97;
output 	ram_block1a121;
output 	ram_block1a145;
output 	ram_block1a169;
output 	ram_block1a49;
output 	ram_block1a73;
output 	ram_block1a1;
output 	ram_block1a25;
output 	ram_block1a98;
output 	ram_block1a122;
output 	ram_block1a146;
output 	ram_block1a170;
output 	ram_block1a50;
output 	ram_block1a74;
output 	ram_block1a2;
output 	ram_block1a26;
output 	ram_block1a99;
output 	ram_block1a123;
output 	ram_block1a147;
output 	ram_block1a171;
output 	ram_block1a51;
output 	ram_block1a75;
output 	ram_block1a3;
output 	ram_block1a27;
output 	ram_block1a100;
output 	ram_block1a124;
output 	ram_block1a148;
output 	ram_block1a172;
output 	ram_block1a52;
output 	ram_block1a76;
output 	ram_block1a4;
output 	ram_block1a28;
output 	ram_block1a101;
output 	ram_block1a125;
output 	ram_block1a149;
output 	ram_block1a173;
output 	ram_block1a53;
output 	ram_block1a77;
output 	ram_block1a5;
output 	ram_block1a29;
output 	ram_block1a102;
output 	ram_block1a126;
output 	ram_block1a150;
output 	ram_block1a174;
output 	ram_block1a54;
output 	ram_block1a78;
output 	ram_block1a6;
output 	ram_block1a30;
output 	ram_block1a103;
output 	ram_block1a127;
output 	ram_block1a151;
output 	ram_block1a175;
output 	ram_block1a55;
output 	ram_block1a79;
output 	ram_block1a7;
output 	ram_block1a31;
output 	ram_block1a104;
output 	ram_block1a128;
output 	ram_block1a152;
output 	ram_block1a176;
output 	ram_block1a56;
output 	ram_block1a80;
output 	ram_block1a8;
output 	ram_block1a32;
output 	ram_block1a105;
output 	ram_block1a129;
output 	ram_block1a153;
output 	ram_block1a177;
output 	ram_block1a57;
output 	ram_block1a81;
output 	ram_block1a9;
output 	ram_block1a33;
output 	ram_block1a106;
output 	ram_block1a130;
output 	ram_block1a154;
output 	ram_block1a178;
output 	ram_block1a58;
output 	ram_block1a82;
output 	ram_block1a10;
output 	ram_block1a34;
output 	ram_block1a107;
output 	ram_block1a131;
output 	ram_block1a155;
output 	ram_block1a179;
output 	ram_block1a59;
output 	ram_block1a83;
output 	ram_block1a11;
output 	ram_block1a35;
output 	ram_block1a108;
output 	ram_block1a132;
output 	ram_block1a156;
output 	ram_block1a180;
output 	ram_block1a60;
output 	ram_block1a84;
output 	ram_block1a12;
output 	ram_block1a36;
output 	ram_block1a109;
output 	ram_block1a133;
output 	ram_block1a157;
output 	ram_block1a181;
output 	ram_block1a61;
output 	ram_block1a85;
output 	ram_block1a13;
output 	ram_block1a37;
output 	ram_block1a110;
output 	ram_block1a134;
output 	ram_block1a158;
output 	ram_block1a182;
output 	ram_block1a62;
output 	ram_block1a86;
output 	ram_block1a14;
output 	ram_block1a38;
output 	ram_block1a111;
output 	ram_block1a135;
output 	ram_block1a159;
output 	ram_block1a183;
output 	ram_block1a63;
output 	ram_block1a87;
output 	ram_block1a15;
output 	ram_block1a39;
output 	ram_block1a112;
output 	ram_block1a136;
output 	ram_block1a160;
output 	ram_block1a184;
output 	ram_block1a64;
output 	ram_block1a88;
output 	ram_block1a16;
output 	ram_block1a40;
output 	ram_block1a113;
output 	ram_block1a137;
output 	ram_block1a161;
output 	ram_block1a185;
output 	ram_block1a65;
output 	ram_block1a89;
output 	ram_block1a17;
output 	ram_block1a41;
output 	ram_block1a114;
output 	ram_block1a138;
output 	ram_block1a162;
output 	ram_block1a186;
output 	ram_block1a66;
output 	ram_block1a90;
output 	ram_block1a18;
output 	ram_block1a42;
output 	ram_block1a115;
output 	ram_block1a139;
output 	ram_block1a163;
output 	ram_block1a187;
output 	ram_block1a67;
output 	ram_block1a91;
output 	ram_block1a19;
output 	ram_block1a43;
output 	ram_block1a116;
output 	ram_block1a140;
output 	ram_block1a164;
output 	ram_block1a188;
output 	ram_block1a68;
output 	ram_block1a92;
output 	ram_block1a20;
output 	ram_block1a44;
output 	ram_block1a117;
output 	ram_block1a141;
output 	ram_block1a165;
output 	ram_block1a189;
output 	ram_block1a69;
output 	ram_block1a93;
output 	ram_block1a21;
output 	ram_block1a45;
output 	ram_block1a118;
output 	ram_block1a142;
output 	ram_block1a166;
output 	ram_block1a190;
output 	ram_block1a70;
output 	ram_block1a94;
output 	ram_block1a22;
output 	ram_block1a46;
output 	ram_block1a119;
output 	ram_block1a143;
output 	ram_block1a167;
output 	ram_block1a191;
output 	ram_block1a71;
output 	ram_block1a95;
output 	ram_block1a23;
output 	ram_block1a47;
input 	[15:0] address_a;
output 	out_address_reg_a_2;
output 	out_address_reg_a_0;
output 	out_address_reg_a_1;
input 	clock0;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_altsyncram_jtf1 auto_generated(
	.ram_block1a961(ram_block1a96),
	.ram_block1a1201(ram_block1a120),
	.ram_block1a1441(ram_block1a144),
	.ram_block1a1681(ram_block1a168),
	.ram_block1a481(ram_block1a48),
	.ram_block1a721(ram_block1a72),
	.ram_block1a01(ram_block1a0),
	.ram_block1a241(ram_block1a24),
	.ram_block1a971(ram_block1a97),
	.ram_block1a1211(ram_block1a121),
	.ram_block1a1451(ram_block1a145),
	.ram_block1a1691(ram_block1a169),
	.ram_block1a491(ram_block1a49),
	.ram_block1a731(ram_block1a73),
	.ram_block1a192(ram_block1a1),
	.ram_block1a251(ram_block1a25),
	.ram_block1a981(ram_block1a98),
	.ram_block1a1221(ram_block1a122),
	.ram_block1a1461(ram_block1a146),
	.ram_block1a1701(ram_block1a170),
	.ram_block1a501(ram_block1a50),
	.ram_block1a741(ram_block1a74),
	.ram_block1a210(ram_block1a2),
	.ram_block1a261(ram_block1a26),
	.ram_block1a991(ram_block1a99),
	.ram_block1a1231(ram_block1a123),
	.ram_block1a1471(ram_block1a147),
	.ram_block1a1711(ram_block1a171),
	.ram_block1a511(ram_block1a51),
	.ram_block1a751(ram_block1a75),
	.ram_block1a310(ram_block1a3),
	.ram_block1a271(ram_block1a27),
	.ram_block1a1001(ram_block1a100),
	.ram_block1a1241(ram_block1a124),
	.ram_block1a1481(ram_block1a148),
	.ram_block1a1721(ram_block1a172),
	.ram_block1a521(ram_block1a52),
	.ram_block1a761(ram_block1a76),
	.ram_block1a410(ram_block1a4),
	.ram_block1a281(ram_block1a28),
	.ram_block1a1011(ram_block1a101),
	.ram_block1a1251(ram_block1a125),
	.ram_block1a1491(ram_block1a149),
	.ram_block1a1731(ram_block1a173),
	.ram_block1a531(ram_block1a53),
	.ram_block1a771(ram_block1a77),
	.ram_block1a510(ram_block1a5),
	.ram_block1a291(ram_block1a29),
	.ram_block1a1021(ram_block1a102),
	.ram_block1a1261(ram_block1a126),
	.ram_block1a1501(ram_block1a150),
	.ram_block1a1741(ram_block1a174),
	.ram_block1a541(ram_block1a54),
	.ram_block1a781(ram_block1a78),
	.ram_block1a610(ram_block1a6),
	.ram_block1a301(ram_block1a30),
	.ram_block1a1031(ram_block1a103),
	.ram_block1a1271(ram_block1a127),
	.ram_block1a1511(ram_block1a151),
	.ram_block1a1751(ram_block1a175),
	.ram_block1a551(ram_block1a55),
	.ram_block1a791(ram_block1a79),
	.ram_block1a710(ram_block1a7),
	.ram_block1a311(ram_block1a31),
	.ram_block1a1041(ram_block1a104),
	.ram_block1a1281(ram_block1a128),
	.ram_block1a1521(ram_block1a152),
	.ram_block1a1761(ram_block1a176),
	.ram_block1a561(ram_block1a56),
	.ram_block1a801(ram_block1a80),
	.ram_block1a810(ram_block1a8),
	.ram_block1a321(ram_block1a32),
	.ram_block1a1051(ram_block1a105),
	.ram_block1a1291(ram_block1a129),
	.ram_block1a1531(ram_block1a153),
	.ram_block1a1771(ram_block1a177),
	.ram_block1a571(ram_block1a57),
	.ram_block1a811(ram_block1a81),
	.ram_block1a910(ram_block1a9),
	.ram_block1a331(ram_block1a33),
	.ram_block1a1061(ram_block1a106),
	.ram_block1a1301(ram_block1a130),
	.ram_block1a1541(ram_block1a154),
	.ram_block1a1781(ram_block1a178),
	.ram_block1a581(ram_block1a58),
	.ram_block1a821(ram_block1a82),
	.ram_block1a1010(ram_block1a10),
	.ram_block1a341(ram_block1a34),
	.ram_block1a1071(ram_block1a107),
	.ram_block1a1311(ram_block1a131),
	.ram_block1a1551(ram_block1a155),
	.ram_block1a1791(ram_block1a179),
	.ram_block1a591(ram_block1a59),
	.ram_block1a831(ram_block1a83),
	.ram_block1a1110(ram_block1a11),
	.ram_block1a351(ram_block1a35),
	.ram_block1a1081(ram_block1a108),
	.ram_block1a1321(ram_block1a132),
	.ram_block1a1561(ram_block1a156),
	.ram_block1a1801(ram_block1a180),
	.ram_block1a601(ram_block1a60),
	.ram_block1a841(ram_block1a84),
	.ram_block1a1210(ram_block1a12),
	.ram_block1a361(ram_block1a36),
	.ram_block1a1091(ram_block1a109),
	.ram_block1a1331(ram_block1a133),
	.ram_block1a1571(ram_block1a157),
	.ram_block1a1811(ram_block1a181),
	.ram_block1a611(ram_block1a61),
	.ram_block1a851(ram_block1a85),
	.ram_block1a1310(ram_block1a13),
	.ram_block1a371(ram_block1a37),
	.ram_block1a1101(ram_block1a110),
	.ram_block1a1341(ram_block1a134),
	.ram_block1a1581(ram_block1a158),
	.ram_block1a1821(ram_block1a182),
	.ram_block1a621(ram_block1a62),
	.ram_block1a861(ram_block1a86),
	.ram_block1a1410(ram_block1a14),
	.ram_block1a381(ram_block1a38),
	.ram_block1a1111(ram_block1a111),
	.ram_block1a1351(ram_block1a135),
	.ram_block1a1591(ram_block1a159),
	.ram_block1a1831(ram_block1a183),
	.ram_block1a631(ram_block1a63),
	.ram_block1a871(ram_block1a87),
	.ram_block1a1510(ram_block1a15),
	.ram_block1a391(ram_block1a39),
	.ram_block1a1121(ram_block1a112),
	.ram_block1a1361(ram_block1a136),
	.ram_block1a1601(ram_block1a160),
	.ram_block1a1841(ram_block1a184),
	.ram_block1a641(ram_block1a64),
	.ram_block1a881(ram_block1a88),
	.ram_block1a1610(ram_block1a16),
	.ram_block1a401(ram_block1a40),
	.ram_block1a1131(ram_block1a113),
	.ram_block1a1371(ram_block1a137),
	.ram_block1a1611(ram_block1a161),
	.ram_block1a1851(ram_block1a185),
	.ram_block1a651(ram_block1a65),
	.ram_block1a891(ram_block1a89),
	.ram_block1a1710(ram_block1a17),
	.ram_block1a411(ram_block1a41),
	.ram_block1a1141(ram_block1a114),
	.ram_block1a1381(ram_block1a138),
	.ram_block1a1621(ram_block1a162),
	.ram_block1a1861(ram_block1a186),
	.ram_block1a661(ram_block1a66),
	.ram_block1a901(ram_block1a90),
	.ram_block1a1810(ram_block1a18),
	.ram_block1a421(ram_block1a42),
	.ram_block1a1151(ram_block1a115),
	.ram_block1a1391(ram_block1a139),
	.ram_block1a1631(ram_block1a163),
	.ram_block1a1871(ram_block1a187),
	.ram_block1a671(ram_block1a67),
	.ram_block1a911(ram_block1a91),
	.ram_block1a193(ram_block1a19),
	.ram_block1a431(ram_block1a43),
	.ram_block1a1161(ram_block1a116),
	.ram_block1a1401(ram_block1a140),
	.ram_block1a1641(ram_block1a164),
	.ram_block1a1881(ram_block1a188),
	.ram_block1a681(ram_block1a68),
	.ram_block1a921(ram_block1a92),
	.ram_block1a201(ram_block1a20),
	.ram_block1a441(ram_block1a44),
	.ram_block1a1171(ram_block1a117),
	.ram_block1a1411(ram_block1a141),
	.ram_block1a1651(ram_block1a165),
	.ram_block1a1891(ram_block1a189),
	.ram_block1a691(ram_block1a69),
	.ram_block1a931(ram_block1a93),
	.ram_block1a211(ram_block1a21),
	.ram_block1a451(ram_block1a45),
	.ram_block1a1181(ram_block1a118),
	.ram_block1a1421(ram_block1a142),
	.ram_block1a1661(ram_block1a166),
	.ram_block1a1901(ram_block1a190),
	.ram_block1a701(ram_block1a70),
	.ram_block1a941(ram_block1a94),
	.ram_block1a221(ram_block1a22),
	.ram_block1a461(ram_block1a46),
	.ram_block1a1191(ram_block1a119),
	.ram_block1a1431(ram_block1a143),
	.ram_block1a1671(ram_block1a167),
	.ram_block1a1911(ram_block1a191),
	.ram_block1a711(ram_block1a71),
	.ram_block1a951(ram_block1a95),
	.ram_block1a231(ram_block1a23),
	.ram_block1a471(ram_block1a47),
	.address_a({address_a[15],address_a[14],address_a[13],address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.out_address_reg_a_2(out_address_reg_a_2),
	.out_address_reg_a_0(out_address_reg_a_0),
	.out_address_reg_a_1(out_address_reg_a_1),
	.clock0(clock0),
	.clocken0(clocken0));

endmodule

module sine_altsyncram_jtf1 (
	ram_block1a961,
	ram_block1a1201,
	ram_block1a1441,
	ram_block1a1681,
	ram_block1a481,
	ram_block1a721,
	ram_block1a01,
	ram_block1a241,
	ram_block1a971,
	ram_block1a1211,
	ram_block1a1451,
	ram_block1a1691,
	ram_block1a491,
	ram_block1a731,
	ram_block1a192,
	ram_block1a251,
	ram_block1a981,
	ram_block1a1221,
	ram_block1a1461,
	ram_block1a1701,
	ram_block1a501,
	ram_block1a741,
	ram_block1a210,
	ram_block1a261,
	ram_block1a991,
	ram_block1a1231,
	ram_block1a1471,
	ram_block1a1711,
	ram_block1a511,
	ram_block1a751,
	ram_block1a310,
	ram_block1a271,
	ram_block1a1001,
	ram_block1a1241,
	ram_block1a1481,
	ram_block1a1721,
	ram_block1a521,
	ram_block1a761,
	ram_block1a410,
	ram_block1a281,
	ram_block1a1011,
	ram_block1a1251,
	ram_block1a1491,
	ram_block1a1731,
	ram_block1a531,
	ram_block1a771,
	ram_block1a510,
	ram_block1a291,
	ram_block1a1021,
	ram_block1a1261,
	ram_block1a1501,
	ram_block1a1741,
	ram_block1a541,
	ram_block1a781,
	ram_block1a610,
	ram_block1a301,
	ram_block1a1031,
	ram_block1a1271,
	ram_block1a1511,
	ram_block1a1751,
	ram_block1a551,
	ram_block1a791,
	ram_block1a710,
	ram_block1a311,
	ram_block1a1041,
	ram_block1a1281,
	ram_block1a1521,
	ram_block1a1761,
	ram_block1a561,
	ram_block1a801,
	ram_block1a810,
	ram_block1a321,
	ram_block1a1051,
	ram_block1a1291,
	ram_block1a1531,
	ram_block1a1771,
	ram_block1a571,
	ram_block1a811,
	ram_block1a910,
	ram_block1a331,
	ram_block1a1061,
	ram_block1a1301,
	ram_block1a1541,
	ram_block1a1781,
	ram_block1a581,
	ram_block1a821,
	ram_block1a1010,
	ram_block1a341,
	ram_block1a1071,
	ram_block1a1311,
	ram_block1a1551,
	ram_block1a1791,
	ram_block1a591,
	ram_block1a831,
	ram_block1a1110,
	ram_block1a351,
	ram_block1a1081,
	ram_block1a1321,
	ram_block1a1561,
	ram_block1a1801,
	ram_block1a601,
	ram_block1a841,
	ram_block1a1210,
	ram_block1a361,
	ram_block1a1091,
	ram_block1a1331,
	ram_block1a1571,
	ram_block1a1811,
	ram_block1a611,
	ram_block1a851,
	ram_block1a1310,
	ram_block1a371,
	ram_block1a1101,
	ram_block1a1341,
	ram_block1a1581,
	ram_block1a1821,
	ram_block1a621,
	ram_block1a861,
	ram_block1a1410,
	ram_block1a381,
	ram_block1a1111,
	ram_block1a1351,
	ram_block1a1591,
	ram_block1a1831,
	ram_block1a631,
	ram_block1a871,
	ram_block1a1510,
	ram_block1a391,
	ram_block1a1121,
	ram_block1a1361,
	ram_block1a1601,
	ram_block1a1841,
	ram_block1a641,
	ram_block1a881,
	ram_block1a1610,
	ram_block1a401,
	ram_block1a1131,
	ram_block1a1371,
	ram_block1a1611,
	ram_block1a1851,
	ram_block1a651,
	ram_block1a891,
	ram_block1a1710,
	ram_block1a411,
	ram_block1a1141,
	ram_block1a1381,
	ram_block1a1621,
	ram_block1a1861,
	ram_block1a661,
	ram_block1a901,
	ram_block1a1810,
	ram_block1a421,
	ram_block1a1151,
	ram_block1a1391,
	ram_block1a1631,
	ram_block1a1871,
	ram_block1a671,
	ram_block1a911,
	ram_block1a193,
	ram_block1a431,
	ram_block1a1161,
	ram_block1a1401,
	ram_block1a1641,
	ram_block1a1881,
	ram_block1a681,
	ram_block1a921,
	ram_block1a201,
	ram_block1a441,
	ram_block1a1171,
	ram_block1a1411,
	ram_block1a1651,
	ram_block1a1891,
	ram_block1a691,
	ram_block1a931,
	ram_block1a211,
	ram_block1a451,
	ram_block1a1181,
	ram_block1a1421,
	ram_block1a1661,
	ram_block1a1901,
	ram_block1a701,
	ram_block1a941,
	ram_block1a221,
	ram_block1a461,
	ram_block1a1191,
	ram_block1a1431,
	ram_block1a1671,
	ram_block1a1911,
	ram_block1a711,
	ram_block1a951,
	ram_block1a231,
	ram_block1a471,
	address_a,
	out_address_reg_a_2,
	out_address_reg_a_0,
	out_address_reg_a_1,
	clock0,
	clocken0)/* synthesis synthesis_greybox=1 */;
output 	ram_block1a961;
output 	ram_block1a1201;
output 	ram_block1a1441;
output 	ram_block1a1681;
output 	ram_block1a481;
output 	ram_block1a721;
output 	ram_block1a01;
output 	ram_block1a241;
output 	ram_block1a971;
output 	ram_block1a1211;
output 	ram_block1a1451;
output 	ram_block1a1691;
output 	ram_block1a491;
output 	ram_block1a731;
output 	ram_block1a192;
output 	ram_block1a251;
output 	ram_block1a981;
output 	ram_block1a1221;
output 	ram_block1a1461;
output 	ram_block1a1701;
output 	ram_block1a501;
output 	ram_block1a741;
output 	ram_block1a210;
output 	ram_block1a261;
output 	ram_block1a991;
output 	ram_block1a1231;
output 	ram_block1a1471;
output 	ram_block1a1711;
output 	ram_block1a511;
output 	ram_block1a751;
output 	ram_block1a310;
output 	ram_block1a271;
output 	ram_block1a1001;
output 	ram_block1a1241;
output 	ram_block1a1481;
output 	ram_block1a1721;
output 	ram_block1a521;
output 	ram_block1a761;
output 	ram_block1a410;
output 	ram_block1a281;
output 	ram_block1a1011;
output 	ram_block1a1251;
output 	ram_block1a1491;
output 	ram_block1a1731;
output 	ram_block1a531;
output 	ram_block1a771;
output 	ram_block1a510;
output 	ram_block1a291;
output 	ram_block1a1021;
output 	ram_block1a1261;
output 	ram_block1a1501;
output 	ram_block1a1741;
output 	ram_block1a541;
output 	ram_block1a781;
output 	ram_block1a610;
output 	ram_block1a301;
output 	ram_block1a1031;
output 	ram_block1a1271;
output 	ram_block1a1511;
output 	ram_block1a1751;
output 	ram_block1a551;
output 	ram_block1a791;
output 	ram_block1a710;
output 	ram_block1a311;
output 	ram_block1a1041;
output 	ram_block1a1281;
output 	ram_block1a1521;
output 	ram_block1a1761;
output 	ram_block1a561;
output 	ram_block1a801;
output 	ram_block1a810;
output 	ram_block1a321;
output 	ram_block1a1051;
output 	ram_block1a1291;
output 	ram_block1a1531;
output 	ram_block1a1771;
output 	ram_block1a571;
output 	ram_block1a811;
output 	ram_block1a910;
output 	ram_block1a331;
output 	ram_block1a1061;
output 	ram_block1a1301;
output 	ram_block1a1541;
output 	ram_block1a1781;
output 	ram_block1a581;
output 	ram_block1a821;
output 	ram_block1a1010;
output 	ram_block1a341;
output 	ram_block1a1071;
output 	ram_block1a1311;
output 	ram_block1a1551;
output 	ram_block1a1791;
output 	ram_block1a591;
output 	ram_block1a831;
output 	ram_block1a1110;
output 	ram_block1a351;
output 	ram_block1a1081;
output 	ram_block1a1321;
output 	ram_block1a1561;
output 	ram_block1a1801;
output 	ram_block1a601;
output 	ram_block1a841;
output 	ram_block1a1210;
output 	ram_block1a361;
output 	ram_block1a1091;
output 	ram_block1a1331;
output 	ram_block1a1571;
output 	ram_block1a1811;
output 	ram_block1a611;
output 	ram_block1a851;
output 	ram_block1a1310;
output 	ram_block1a371;
output 	ram_block1a1101;
output 	ram_block1a1341;
output 	ram_block1a1581;
output 	ram_block1a1821;
output 	ram_block1a621;
output 	ram_block1a861;
output 	ram_block1a1410;
output 	ram_block1a381;
output 	ram_block1a1111;
output 	ram_block1a1351;
output 	ram_block1a1591;
output 	ram_block1a1831;
output 	ram_block1a631;
output 	ram_block1a871;
output 	ram_block1a1510;
output 	ram_block1a391;
output 	ram_block1a1121;
output 	ram_block1a1361;
output 	ram_block1a1601;
output 	ram_block1a1841;
output 	ram_block1a641;
output 	ram_block1a881;
output 	ram_block1a1610;
output 	ram_block1a401;
output 	ram_block1a1131;
output 	ram_block1a1371;
output 	ram_block1a1611;
output 	ram_block1a1851;
output 	ram_block1a651;
output 	ram_block1a891;
output 	ram_block1a1710;
output 	ram_block1a411;
output 	ram_block1a1141;
output 	ram_block1a1381;
output 	ram_block1a1621;
output 	ram_block1a1861;
output 	ram_block1a661;
output 	ram_block1a901;
output 	ram_block1a1810;
output 	ram_block1a421;
output 	ram_block1a1151;
output 	ram_block1a1391;
output 	ram_block1a1631;
output 	ram_block1a1871;
output 	ram_block1a671;
output 	ram_block1a911;
output 	ram_block1a193;
output 	ram_block1a431;
output 	ram_block1a1161;
output 	ram_block1a1401;
output 	ram_block1a1641;
output 	ram_block1a1881;
output 	ram_block1a681;
output 	ram_block1a921;
output 	ram_block1a201;
output 	ram_block1a441;
output 	ram_block1a1171;
output 	ram_block1a1411;
output 	ram_block1a1651;
output 	ram_block1a1891;
output 	ram_block1a691;
output 	ram_block1a931;
output 	ram_block1a211;
output 	ram_block1a451;
output 	ram_block1a1181;
output 	ram_block1a1421;
output 	ram_block1a1661;
output 	ram_block1a1901;
output 	ram_block1a701;
output 	ram_block1a941;
output 	ram_block1a221;
output 	ram_block1a461;
output 	ram_block1a1191;
output 	ram_block1a1431;
output 	ram_block1a1671;
output 	ram_block1a1911;
output 	ram_block1a711;
output 	ram_block1a951;
output 	ram_block1a231;
output 	ram_block1a471;
input 	[15:0] address_a;
output 	out_address_reg_a_2;
output 	out_address_reg_a_0;
output 	out_address_reg_a_1;
input 	clock0;
input 	clocken0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \address_reg_a[2]~q ;
wire \address_reg_a[0]~q ;
wire \address_reg_a[1]~q ;

wire [143:0] ram_block1a96_PORTADATAOUT_bus;
wire [143:0] ram_block1a120_PORTADATAOUT_bus;
wire [143:0] ram_block1a144_PORTADATAOUT_bus;
wire [143:0] ram_block1a168_PORTADATAOUT_bus;
wire [143:0] ram_block1a48_PORTADATAOUT_bus;
wire [143:0] ram_block1a72_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a97_PORTADATAOUT_bus;
wire [143:0] ram_block1a121_PORTADATAOUT_bus;
wire [143:0] ram_block1a145_PORTADATAOUT_bus;
wire [143:0] ram_block1a169_PORTADATAOUT_bus;
wire [143:0] ram_block1a49_PORTADATAOUT_bus;
wire [143:0] ram_block1a73_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a98_PORTADATAOUT_bus;
wire [143:0] ram_block1a122_PORTADATAOUT_bus;
wire [143:0] ram_block1a146_PORTADATAOUT_bus;
wire [143:0] ram_block1a170_PORTADATAOUT_bus;
wire [143:0] ram_block1a50_PORTADATAOUT_bus;
wire [143:0] ram_block1a74_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a99_PORTADATAOUT_bus;
wire [143:0] ram_block1a123_PORTADATAOUT_bus;
wire [143:0] ram_block1a147_PORTADATAOUT_bus;
wire [143:0] ram_block1a171_PORTADATAOUT_bus;
wire [143:0] ram_block1a51_PORTADATAOUT_bus;
wire [143:0] ram_block1a75_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a100_PORTADATAOUT_bus;
wire [143:0] ram_block1a124_PORTADATAOUT_bus;
wire [143:0] ram_block1a148_PORTADATAOUT_bus;
wire [143:0] ram_block1a172_PORTADATAOUT_bus;
wire [143:0] ram_block1a52_PORTADATAOUT_bus;
wire [143:0] ram_block1a76_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a101_PORTADATAOUT_bus;
wire [143:0] ram_block1a125_PORTADATAOUT_bus;
wire [143:0] ram_block1a149_PORTADATAOUT_bus;
wire [143:0] ram_block1a173_PORTADATAOUT_bus;
wire [143:0] ram_block1a53_PORTADATAOUT_bus;
wire [143:0] ram_block1a77_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a102_PORTADATAOUT_bus;
wire [143:0] ram_block1a126_PORTADATAOUT_bus;
wire [143:0] ram_block1a150_PORTADATAOUT_bus;
wire [143:0] ram_block1a174_PORTADATAOUT_bus;
wire [143:0] ram_block1a54_PORTADATAOUT_bus;
wire [143:0] ram_block1a78_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a103_PORTADATAOUT_bus;
wire [143:0] ram_block1a127_PORTADATAOUT_bus;
wire [143:0] ram_block1a151_PORTADATAOUT_bus;
wire [143:0] ram_block1a175_PORTADATAOUT_bus;
wire [143:0] ram_block1a55_PORTADATAOUT_bus;
wire [143:0] ram_block1a79_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a104_PORTADATAOUT_bus;
wire [143:0] ram_block1a128_PORTADATAOUT_bus;
wire [143:0] ram_block1a152_PORTADATAOUT_bus;
wire [143:0] ram_block1a176_PORTADATAOUT_bus;
wire [143:0] ram_block1a56_PORTADATAOUT_bus;
wire [143:0] ram_block1a80_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a32_PORTADATAOUT_bus;
wire [143:0] ram_block1a105_PORTADATAOUT_bus;
wire [143:0] ram_block1a129_PORTADATAOUT_bus;
wire [143:0] ram_block1a153_PORTADATAOUT_bus;
wire [143:0] ram_block1a177_PORTADATAOUT_bus;
wire [143:0] ram_block1a57_PORTADATAOUT_bus;
wire [143:0] ram_block1a81_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a33_PORTADATAOUT_bus;
wire [143:0] ram_block1a106_PORTADATAOUT_bus;
wire [143:0] ram_block1a130_PORTADATAOUT_bus;
wire [143:0] ram_block1a154_PORTADATAOUT_bus;
wire [143:0] ram_block1a178_PORTADATAOUT_bus;
wire [143:0] ram_block1a58_PORTADATAOUT_bus;
wire [143:0] ram_block1a82_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a34_PORTADATAOUT_bus;
wire [143:0] ram_block1a107_PORTADATAOUT_bus;
wire [143:0] ram_block1a131_PORTADATAOUT_bus;
wire [143:0] ram_block1a155_PORTADATAOUT_bus;
wire [143:0] ram_block1a179_PORTADATAOUT_bus;
wire [143:0] ram_block1a59_PORTADATAOUT_bus;
wire [143:0] ram_block1a83_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a35_PORTADATAOUT_bus;
wire [143:0] ram_block1a108_PORTADATAOUT_bus;
wire [143:0] ram_block1a132_PORTADATAOUT_bus;
wire [143:0] ram_block1a156_PORTADATAOUT_bus;
wire [143:0] ram_block1a180_PORTADATAOUT_bus;
wire [143:0] ram_block1a60_PORTADATAOUT_bus;
wire [143:0] ram_block1a84_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a36_PORTADATAOUT_bus;
wire [143:0] ram_block1a109_PORTADATAOUT_bus;
wire [143:0] ram_block1a133_PORTADATAOUT_bus;
wire [143:0] ram_block1a157_PORTADATAOUT_bus;
wire [143:0] ram_block1a181_PORTADATAOUT_bus;
wire [143:0] ram_block1a61_PORTADATAOUT_bus;
wire [143:0] ram_block1a85_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a37_PORTADATAOUT_bus;
wire [143:0] ram_block1a110_PORTADATAOUT_bus;
wire [143:0] ram_block1a134_PORTADATAOUT_bus;
wire [143:0] ram_block1a158_PORTADATAOUT_bus;
wire [143:0] ram_block1a182_PORTADATAOUT_bus;
wire [143:0] ram_block1a62_PORTADATAOUT_bus;
wire [143:0] ram_block1a86_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a38_PORTADATAOUT_bus;
wire [143:0] ram_block1a111_PORTADATAOUT_bus;
wire [143:0] ram_block1a135_PORTADATAOUT_bus;
wire [143:0] ram_block1a159_PORTADATAOUT_bus;
wire [143:0] ram_block1a183_PORTADATAOUT_bus;
wire [143:0] ram_block1a63_PORTADATAOUT_bus;
wire [143:0] ram_block1a87_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a39_PORTADATAOUT_bus;
wire [143:0] ram_block1a112_PORTADATAOUT_bus;
wire [143:0] ram_block1a136_PORTADATAOUT_bus;
wire [143:0] ram_block1a160_PORTADATAOUT_bus;
wire [143:0] ram_block1a184_PORTADATAOUT_bus;
wire [143:0] ram_block1a64_PORTADATAOUT_bus;
wire [143:0] ram_block1a88_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a40_PORTADATAOUT_bus;
wire [143:0] ram_block1a113_PORTADATAOUT_bus;
wire [143:0] ram_block1a137_PORTADATAOUT_bus;
wire [143:0] ram_block1a161_PORTADATAOUT_bus;
wire [143:0] ram_block1a185_PORTADATAOUT_bus;
wire [143:0] ram_block1a65_PORTADATAOUT_bus;
wire [143:0] ram_block1a89_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a41_PORTADATAOUT_bus;
wire [143:0] ram_block1a114_PORTADATAOUT_bus;
wire [143:0] ram_block1a138_PORTADATAOUT_bus;
wire [143:0] ram_block1a162_PORTADATAOUT_bus;
wire [143:0] ram_block1a186_PORTADATAOUT_bus;
wire [143:0] ram_block1a66_PORTADATAOUT_bus;
wire [143:0] ram_block1a90_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a42_PORTADATAOUT_bus;
wire [143:0] ram_block1a115_PORTADATAOUT_bus;
wire [143:0] ram_block1a139_PORTADATAOUT_bus;
wire [143:0] ram_block1a163_PORTADATAOUT_bus;
wire [143:0] ram_block1a187_PORTADATAOUT_bus;
wire [143:0] ram_block1a67_PORTADATAOUT_bus;
wire [143:0] ram_block1a91_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a43_PORTADATAOUT_bus;
wire [143:0] ram_block1a116_PORTADATAOUT_bus;
wire [143:0] ram_block1a140_PORTADATAOUT_bus;
wire [143:0] ram_block1a164_PORTADATAOUT_bus;
wire [143:0] ram_block1a188_PORTADATAOUT_bus;
wire [143:0] ram_block1a68_PORTADATAOUT_bus;
wire [143:0] ram_block1a92_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a44_PORTADATAOUT_bus;
wire [143:0] ram_block1a117_PORTADATAOUT_bus;
wire [143:0] ram_block1a141_PORTADATAOUT_bus;
wire [143:0] ram_block1a165_PORTADATAOUT_bus;
wire [143:0] ram_block1a189_PORTADATAOUT_bus;
wire [143:0] ram_block1a69_PORTADATAOUT_bus;
wire [143:0] ram_block1a93_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a45_PORTADATAOUT_bus;
wire [143:0] ram_block1a118_PORTADATAOUT_bus;
wire [143:0] ram_block1a142_PORTADATAOUT_bus;
wire [143:0] ram_block1a166_PORTADATAOUT_bus;
wire [143:0] ram_block1a190_PORTADATAOUT_bus;
wire [143:0] ram_block1a70_PORTADATAOUT_bus;
wire [143:0] ram_block1a94_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a46_PORTADATAOUT_bus;
wire [143:0] ram_block1a119_PORTADATAOUT_bus;
wire [143:0] ram_block1a143_PORTADATAOUT_bus;
wire [143:0] ram_block1a167_PORTADATAOUT_bus;
wire [143:0] ram_block1a191_PORTADATAOUT_bus;
wire [143:0] ram_block1a71_PORTADATAOUT_bus;
wire [143:0] ram_block1a95_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a47_PORTADATAOUT_bus;

assign ram_block1a961 = ram_block1a96_PORTADATAOUT_bus[0];

assign ram_block1a1201 = ram_block1a120_PORTADATAOUT_bus[0];

assign ram_block1a1441 = ram_block1a144_PORTADATAOUT_bus[0];

assign ram_block1a1681 = ram_block1a168_PORTADATAOUT_bus[0];

assign ram_block1a481 = ram_block1a48_PORTADATAOUT_bus[0];

assign ram_block1a721 = ram_block1a72_PORTADATAOUT_bus[0];

assign ram_block1a01 = ram_block1a0_PORTADATAOUT_bus[0];

assign ram_block1a241 = ram_block1a24_PORTADATAOUT_bus[0];

assign ram_block1a971 = ram_block1a97_PORTADATAOUT_bus[0];

assign ram_block1a1211 = ram_block1a121_PORTADATAOUT_bus[0];

assign ram_block1a1451 = ram_block1a145_PORTADATAOUT_bus[0];

assign ram_block1a1691 = ram_block1a169_PORTADATAOUT_bus[0];

assign ram_block1a491 = ram_block1a49_PORTADATAOUT_bus[0];

assign ram_block1a731 = ram_block1a73_PORTADATAOUT_bus[0];

assign ram_block1a192 = ram_block1a1_PORTADATAOUT_bus[0];

assign ram_block1a251 = ram_block1a25_PORTADATAOUT_bus[0];

assign ram_block1a981 = ram_block1a98_PORTADATAOUT_bus[0];

assign ram_block1a1221 = ram_block1a122_PORTADATAOUT_bus[0];

assign ram_block1a1461 = ram_block1a146_PORTADATAOUT_bus[0];

assign ram_block1a1701 = ram_block1a170_PORTADATAOUT_bus[0];

assign ram_block1a501 = ram_block1a50_PORTADATAOUT_bus[0];

assign ram_block1a741 = ram_block1a74_PORTADATAOUT_bus[0];

assign ram_block1a210 = ram_block1a2_PORTADATAOUT_bus[0];

assign ram_block1a261 = ram_block1a26_PORTADATAOUT_bus[0];

assign ram_block1a991 = ram_block1a99_PORTADATAOUT_bus[0];

assign ram_block1a1231 = ram_block1a123_PORTADATAOUT_bus[0];

assign ram_block1a1471 = ram_block1a147_PORTADATAOUT_bus[0];

assign ram_block1a1711 = ram_block1a171_PORTADATAOUT_bus[0];

assign ram_block1a511 = ram_block1a51_PORTADATAOUT_bus[0];

assign ram_block1a751 = ram_block1a75_PORTADATAOUT_bus[0];

assign ram_block1a310 = ram_block1a3_PORTADATAOUT_bus[0];

assign ram_block1a271 = ram_block1a27_PORTADATAOUT_bus[0];

assign ram_block1a1001 = ram_block1a100_PORTADATAOUT_bus[0];

assign ram_block1a1241 = ram_block1a124_PORTADATAOUT_bus[0];

assign ram_block1a1481 = ram_block1a148_PORTADATAOUT_bus[0];

assign ram_block1a1721 = ram_block1a172_PORTADATAOUT_bus[0];

assign ram_block1a521 = ram_block1a52_PORTADATAOUT_bus[0];

assign ram_block1a761 = ram_block1a76_PORTADATAOUT_bus[0];

assign ram_block1a410 = ram_block1a4_PORTADATAOUT_bus[0];

assign ram_block1a281 = ram_block1a28_PORTADATAOUT_bus[0];

assign ram_block1a1011 = ram_block1a101_PORTADATAOUT_bus[0];

assign ram_block1a1251 = ram_block1a125_PORTADATAOUT_bus[0];

assign ram_block1a1491 = ram_block1a149_PORTADATAOUT_bus[0];

assign ram_block1a1731 = ram_block1a173_PORTADATAOUT_bus[0];

assign ram_block1a531 = ram_block1a53_PORTADATAOUT_bus[0];

assign ram_block1a771 = ram_block1a77_PORTADATAOUT_bus[0];

assign ram_block1a510 = ram_block1a5_PORTADATAOUT_bus[0];

assign ram_block1a291 = ram_block1a29_PORTADATAOUT_bus[0];

assign ram_block1a1021 = ram_block1a102_PORTADATAOUT_bus[0];

assign ram_block1a1261 = ram_block1a126_PORTADATAOUT_bus[0];

assign ram_block1a1501 = ram_block1a150_PORTADATAOUT_bus[0];

assign ram_block1a1741 = ram_block1a174_PORTADATAOUT_bus[0];

assign ram_block1a541 = ram_block1a54_PORTADATAOUT_bus[0];

assign ram_block1a781 = ram_block1a78_PORTADATAOUT_bus[0];

assign ram_block1a610 = ram_block1a6_PORTADATAOUT_bus[0];

assign ram_block1a301 = ram_block1a30_PORTADATAOUT_bus[0];

assign ram_block1a1031 = ram_block1a103_PORTADATAOUT_bus[0];

assign ram_block1a1271 = ram_block1a127_PORTADATAOUT_bus[0];

assign ram_block1a1511 = ram_block1a151_PORTADATAOUT_bus[0];

assign ram_block1a1751 = ram_block1a175_PORTADATAOUT_bus[0];

assign ram_block1a551 = ram_block1a55_PORTADATAOUT_bus[0];

assign ram_block1a791 = ram_block1a79_PORTADATAOUT_bus[0];

assign ram_block1a710 = ram_block1a7_PORTADATAOUT_bus[0];

assign ram_block1a311 = ram_block1a31_PORTADATAOUT_bus[0];

assign ram_block1a1041 = ram_block1a104_PORTADATAOUT_bus[0];

assign ram_block1a1281 = ram_block1a128_PORTADATAOUT_bus[0];

assign ram_block1a1521 = ram_block1a152_PORTADATAOUT_bus[0];

assign ram_block1a1761 = ram_block1a176_PORTADATAOUT_bus[0];

assign ram_block1a561 = ram_block1a56_PORTADATAOUT_bus[0];

assign ram_block1a801 = ram_block1a80_PORTADATAOUT_bus[0];

assign ram_block1a810 = ram_block1a8_PORTADATAOUT_bus[0];

assign ram_block1a321 = ram_block1a32_PORTADATAOUT_bus[0];

assign ram_block1a1051 = ram_block1a105_PORTADATAOUT_bus[0];

assign ram_block1a1291 = ram_block1a129_PORTADATAOUT_bus[0];

assign ram_block1a1531 = ram_block1a153_PORTADATAOUT_bus[0];

assign ram_block1a1771 = ram_block1a177_PORTADATAOUT_bus[0];

assign ram_block1a571 = ram_block1a57_PORTADATAOUT_bus[0];

assign ram_block1a811 = ram_block1a81_PORTADATAOUT_bus[0];

assign ram_block1a910 = ram_block1a9_PORTADATAOUT_bus[0];

assign ram_block1a331 = ram_block1a33_PORTADATAOUT_bus[0];

assign ram_block1a1061 = ram_block1a106_PORTADATAOUT_bus[0];

assign ram_block1a1301 = ram_block1a130_PORTADATAOUT_bus[0];

assign ram_block1a1541 = ram_block1a154_PORTADATAOUT_bus[0];

assign ram_block1a1781 = ram_block1a178_PORTADATAOUT_bus[0];

assign ram_block1a581 = ram_block1a58_PORTADATAOUT_bus[0];

assign ram_block1a821 = ram_block1a82_PORTADATAOUT_bus[0];

assign ram_block1a1010 = ram_block1a10_PORTADATAOUT_bus[0];

assign ram_block1a341 = ram_block1a34_PORTADATAOUT_bus[0];

assign ram_block1a1071 = ram_block1a107_PORTADATAOUT_bus[0];

assign ram_block1a1311 = ram_block1a131_PORTADATAOUT_bus[0];

assign ram_block1a1551 = ram_block1a155_PORTADATAOUT_bus[0];

assign ram_block1a1791 = ram_block1a179_PORTADATAOUT_bus[0];

assign ram_block1a591 = ram_block1a59_PORTADATAOUT_bus[0];

assign ram_block1a831 = ram_block1a83_PORTADATAOUT_bus[0];

assign ram_block1a1110 = ram_block1a11_PORTADATAOUT_bus[0];

assign ram_block1a351 = ram_block1a35_PORTADATAOUT_bus[0];

assign ram_block1a1081 = ram_block1a108_PORTADATAOUT_bus[0];

assign ram_block1a1321 = ram_block1a132_PORTADATAOUT_bus[0];

assign ram_block1a1561 = ram_block1a156_PORTADATAOUT_bus[0];

assign ram_block1a1801 = ram_block1a180_PORTADATAOUT_bus[0];

assign ram_block1a601 = ram_block1a60_PORTADATAOUT_bus[0];

assign ram_block1a841 = ram_block1a84_PORTADATAOUT_bus[0];

assign ram_block1a1210 = ram_block1a12_PORTADATAOUT_bus[0];

assign ram_block1a361 = ram_block1a36_PORTADATAOUT_bus[0];

assign ram_block1a1091 = ram_block1a109_PORTADATAOUT_bus[0];

assign ram_block1a1331 = ram_block1a133_PORTADATAOUT_bus[0];

assign ram_block1a1571 = ram_block1a157_PORTADATAOUT_bus[0];

assign ram_block1a1811 = ram_block1a181_PORTADATAOUT_bus[0];

assign ram_block1a611 = ram_block1a61_PORTADATAOUT_bus[0];

assign ram_block1a851 = ram_block1a85_PORTADATAOUT_bus[0];

assign ram_block1a1310 = ram_block1a13_PORTADATAOUT_bus[0];

assign ram_block1a371 = ram_block1a37_PORTADATAOUT_bus[0];

assign ram_block1a1101 = ram_block1a110_PORTADATAOUT_bus[0];

assign ram_block1a1341 = ram_block1a134_PORTADATAOUT_bus[0];

assign ram_block1a1581 = ram_block1a158_PORTADATAOUT_bus[0];

assign ram_block1a1821 = ram_block1a182_PORTADATAOUT_bus[0];

assign ram_block1a621 = ram_block1a62_PORTADATAOUT_bus[0];

assign ram_block1a861 = ram_block1a86_PORTADATAOUT_bus[0];

assign ram_block1a1410 = ram_block1a14_PORTADATAOUT_bus[0];

assign ram_block1a381 = ram_block1a38_PORTADATAOUT_bus[0];

assign ram_block1a1111 = ram_block1a111_PORTADATAOUT_bus[0];

assign ram_block1a1351 = ram_block1a135_PORTADATAOUT_bus[0];

assign ram_block1a1591 = ram_block1a159_PORTADATAOUT_bus[0];

assign ram_block1a1831 = ram_block1a183_PORTADATAOUT_bus[0];

assign ram_block1a631 = ram_block1a63_PORTADATAOUT_bus[0];

assign ram_block1a871 = ram_block1a87_PORTADATAOUT_bus[0];

assign ram_block1a1510 = ram_block1a15_PORTADATAOUT_bus[0];

assign ram_block1a391 = ram_block1a39_PORTADATAOUT_bus[0];

assign ram_block1a1121 = ram_block1a112_PORTADATAOUT_bus[0];

assign ram_block1a1361 = ram_block1a136_PORTADATAOUT_bus[0];

assign ram_block1a1601 = ram_block1a160_PORTADATAOUT_bus[0];

assign ram_block1a1841 = ram_block1a184_PORTADATAOUT_bus[0];

assign ram_block1a641 = ram_block1a64_PORTADATAOUT_bus[0];

assign ram_block1a881 = ram_block1a88_PORTADATAOUT_bus[0];

assign ram_block1a1610 = ram_block1a16_PORTADATAOUT_bus[0];

assign ram_block1a401 = ram_block1a40_PORTADATAOUT_bus[0];

assign ram_block1a1131 = ram_block1a113_PORTADATAOUT_bus[0];

assign ram_block1a1371 = ram_block1a137_PORTADATAOUT_bus[0];

assign ram_block1a1611 = ram_block1a161_PORTADATAOUT_bus[0];

assign ram_block1a1851 = ram_block1a185_PORTADATAOUT_bus[0];

assign ram_block1a651 = ram_block1a65_PORTADATAOUT_bus[0];

assign ram_block1a891 = ram_block1a89_PORTADATAOUT_bus[0];

assign ram_block1a1710 = ram_block1a17_PORTADATAOUT_bus[0];

assign ram_block1a411 = ram_block1a41_PORTADATAOUT_bus[0];

assign ram_block1a1141 = ram_block1a114_PORTADATAOUT_bus[0];

assign ram_block1a1381 = ram_block1a138_PORTADATAOUT_bus[0];

assign ram_block1a1621 = ram_block1a162_PORTADATAOUT_bus[0];

assign ram_block1a1861 = ram_block1a186_PORTADATAOUT_bus[0];

assign ram_block1a661 = ram_block1a66_PORTADATAOUT_bus[0];

assign ram_block1a901 = ram_block1a90_PORTADATAOUT_bus[0];

assign ram_block1a1810 = ram_block1a18_PORTADATAOUT_bus[0];

assign ram_block1a421 = ram_block1a42_PORTADATAOUT_bus[0];

assign ram_block1a1151 = ram_block1a115_PORTADATAOUT_bus[0];

assign ram_block1a1391 = ram_block1a139_PORTADATAOUT_bus[0];

assign ram_block1a1631 = ram_block1a163_PORTADATAOUT_bus[0];

assign ram_block1a1871 = ram_block1a187_PORTADATAOUT_bus[0];

assign ram_block1a671 = ram_block1a67_PORTADATAOUT_bus[0];

assign ram_block1a911 = ram_block1a91_PORTADATAOUT_bus[0];

assign ram_block1a193 = ram_block1a19_PORTADATAOUT_bus[0];

assign ram_block1a431 = ram_block1a43_PORTADATAOUT_bus[0];

assign ram_block1a1161 = ram_block1a116_PORTADATAOUT_bus[0];

assign ram_block1a1401 = ram_block1a140_PORTADATAOUT_bus[0];

assign ram_block1a1641 = ram_block1a164_PORTADATAOUT_bus[0];

assign ram_block1a1881 = ram_block1a188_PORTADATAOUT_bus[0];

assign ram_block1a681 = ram_block1a68_PORTADATAOUT_bus[0];

assign ram_block1a921 = ram_block1a92_PORTADATAOUT_bus[0];

assign ram_block1a201 = ram_block1a20_PORTADATAOUT_bus[0];

assign ram_block1a441 = ram_block1a44_PORTADATAOUT_bus[0];

assign ram_block1a1171 = ram_block1a117_PORTADATAOUT_bus[0];

assign ram_block1a1411 = ram_block1a141_PORTADATAOUT_bus[0];

assign ram_block1a1651 = ram_block1a165_PORTADATAOUT_bus[0];

assign ram_block1a1891 = ram_block1a189_PORTADATAOUT_bus[0];

assign ram_block1a691 = ram_block1a69_PORTADATAOUT_bus[0];

assign ram_block1a931 = ram_block1a93_PORTADATAOUT_bus[0];

assign ram_block1a211 = ram_block1a21_PORTADATAOUT_bus[0];

assign ram_block1a451 = ram_block1a45_PORTADATAOUT_bus[0];

assign ram_block1a1181 = ram_block1a118_PORTADATAOUT_bus[0];

assign ram_block1a1421 = ram_block1a142_PORTADATAOUT_bus[0];

assign ram_block1a1661 = ram_block1a166_PORTADATAOUT_bus[0];

assign ram_block1a1901 = ram_block1a190_PORTADATAOUT_bus[0];

assign ram_block1a701 = ram_block1a70_PORTADATAOUT_bus[0];

assign ram_block1a941 = ram_block1a94_PORTADATAOUT_bus[0];

assign ram_block1a221 = ram_block1a22_PORTADATAOUT_bus[0];

assign ram_block1a461 = ram_block1a46_PORTADATAOUT_bus[0];

assign ram_block1a1191 = ram_block1a119_PORTADATAOUT_bus[0];

assign ram_block1a1431 = ram_block1a143_PORTADATAOUT_bus[0];

assign ram_block1a1671 = ram_block1a167_PORTADATAOUT_bus[0];

assign ram_block1a1911 = ram_block1a191_PORTADATAOUT_bus[0];

assign ram_block1a711 = ram_block1a71_PORTADATAOUT_bus[0];

assign ram_block1a951 = ram_block1a95_PORTADATAOUT_bus[0];

assign ram_block1a231 = ram_block1a23_PORTADATAOUT_bus[0];

assign ram_block1a471 = ram_block1a47_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a96(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a96_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a96.clk0_core_clock_enable = "ena0";
defparam ram_block1a96.clk0_input_clock_enable = "ena0";
defparam ram_block1a96.clk0_output_clock_enable = "ena0";
defparam ram_block1a96.data_interleave_offset_in_bits = 1;
defparam ram_block1a96.data_interleave_width_in_bits = 1;
defparam ram_block1a96.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a96.init_file_layout = "port_a";
defparam ram_block1a96.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a96.operation_mode = "rom";
defparam ram_block1a96.port_a_address_clear = "none";
defparam ram_block1a96.port_a_address_width = 13;
defparam ram_block1a96.port_a_data_out_clear = "none";
defparam ram_block1a96.port_a_data_out_clock = "clock0";
defparam ram_block1a96.port_a_data_width = 1;
defparam ram_block1a96.port_a_first_address = 32768;
defparam ram_block1a96.port_a_first_bit_number = 0;
defparam ram_block1a96.port_a_last_address = 40959;
defparam ram_block1a96.port_a_logical_ram_depth = 65536;
defparam ram_block1a96.port_a_logical_ram_width = 24;
defparam ram_block1a96.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a96.ram_block_type = "auto";
defparam ram_block1a96.mem_init3 = "6A5987C3B6A933C1E65A967001C94D6E7FF335549C00734A9670039B55B70FC725549C1C19A5699E03992AD98FF19A5499C03892A931FFC6D296C7FF192AB67001896B49C00392D691800E6D55B3C03CDAAB638079B554CC0019B556C700E36AAD9838392D4B30FE19B55B31FF0C955267C3E64AAD987F0CD2A598FFC66952CC3FC7255533020736AA59C0039B556CC3F866D5491800736AA931FFC76D5499C00E64AAD98FFE32575271FF8CD2AD33800E65AA4987FC7252D64780F1B4A9663FFC66B52D8E00F32D5499C00732554918003994AD263FFC66D55B31FFE334AA49C7FE33294A661FE1C96A9663C1F3B6AADB9F07CEDAAB667C1F1B6AA933800732";
defparam ram_block1a96.mem_init2 = "555263C03CCD2AD263FFE336AAB663FFC725AA591C00399296B661FF8E6D55499E0038DB55699C0C0E64AAA4CC1FC39B4AB49CFC3E334AAB667803CEDAAA933C0038DB554B31F07C66D5549987FC39B4AA5B183F87325556DCF001C64B55A4C7801C6695549987FF0C495B526707E0E64AD29271FFF8E49555B6383C0E669552D9C3FF8E64A56B663C00F39255524CF00038C96AA5B31F83F19B4AAD26707F87336AAADB187FF0E64A54A49C7C07C66D2AAD333C001C66D2AA5938F00F8CC94A94998F003C664A54A49CF00071992A4AD331E003C664A55AD99C7FFC31B2D5569B187FFC3992D554B331F007C664B554B6670FFF0E66DAAA96CCF0FF838C92D5";
defparam ram_block1a96.mem_init1 = "5A498E1FFC1CCDA55569B38F803E39B69554B6671FFFF1CCDA5552DB31E0003C66495554B26383FF0719B6B55292671F003E39925AAA524CE3F007C7336D4A95B6661F001E18D929556B6CC70FFFE1C66DA5554B64E70FFFE1C664B5AAD69331C3FFFC38CDB4AAAA5B6638FF0FE1CE4DAD5552DB338F8001F1CCDB6A96A96CCC70FFFF839CDB6B5552926661E000078E664B5AAAD693338F00E00F18CDB4A555AD26CE70FE01FC798D92D4AAB5A4998C3C000078E3324B5AAA94B6CCC70FC007F1E732692B555A96C99CE1E00007C39CC9B4A5555296D998C780FFF81E399992D2B554AD2D9998E1F00001F0E33336D2B5555A96D9998E3C07FFC078E33326D2";
defparam ram_block1a96.mem_init0 = "9555552D24999CE1E07FFFC0F1C6336496952AA95292C9999C70FC00000FC38C6666DB4A554B556B4926CCE71C3E007F003E1E31999B24B4AD55554AD6D26CCCC638783FF007FE0F0E399C99B6D2D6AD5554AB5A4B64CCCCE30E1F01FFFFFC07C3C718CCCC9B6DA52954AAAA55294B6DB66CCC671870F07F00000003F83E1C71CC66664D924B4B5A955AAAAA556A5292DB6D933667318C71C3C3E07F0007FFC001FE07C3C38718E7339999B364DB6DA4B4A52B56AA5555555552AB54AD6B5A5B4924924D93266CCCCC667318E718E3C70E1E1E1F07C0FC07F803FFC00007FFFFFFF000007FFE007FC01FC07F03F03F07E0F83E0F07C3E1E0F0F0787878787878";

cyclonev_ram_block ram_block1a120(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a120_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a120.clk0_core_clock_enable = "ena0";
defparam ram_block1a120.clk0_input_clock_enable = "ena0";
defparam ram_block1a120.clk0_output_clock_enable = "ena0";
defparam ram_block1a120.data_interleave_offset_in_bits = 1;
defparam ram_block1a120.data_interleave_width_in_bits = 1;
defparam ram_block1a120.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a120.init_file_layout = "port_a";
defparam ram_block1a120.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a120.operation_mode = "rom";
defparam ram_block1a120.port_a_address_clear = "none";
defparam ram_block1a120.port_a_address_width = 13;
defparam ram_block1a120.port_a_data_out_clear = "none";
defparam ram_block1a120.port_a_data_out_clock = "clock0";
defparam ram_block1a120.port_a_data_width = 1;
defparam ram_block1a120.port_a_first_address = 40960;
defparam ram_block1a120.port_a_first_bit_number = 0;
defparam ram_block1a120.port_a_last_address = 49151;
defparam ram_block1a120.port_a_logical_ram_depth = 65536;
defparam ram_block1a120.port_a_logical_ram_width = 24;
defparam ram_block1a120.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a120.ram_block_type = "auto";
defparam ram_block1a120.mem_init3 = "E35563F8954C7C655B003252701DAACFFCDA58FC6D498066A99FE65598066A99FC6D49C1CD34C00DAA67F1A5B3FF2559C1CD54E0392930064ACC01DAB70076ADC01DAB30064A4C0192D380E556E073559E3C9523FE6D6CFF1AA98F8CAB60836ACC0196D380ED567073559E3C9527FF2548FF89523FE2549E3C956707355B80E4A4C00CAA47F9B5270396931E325B38792B63F9956C00C969C072AB701DAA9C0325260065523FC4AB700ED567DE6D6CFF9A4B3FE6D6CF7CD54E01DAACFFCDA58FE25563F8DAD9EF9AA980192D380ED56E0396930832AB38792A67FCCA93C39A69870DA930064A4C00CAACFFCDAD9FF36A4F0F2D6C7F12A91FC6D49C0E6AB3C79A";
defparam ram_block1a120.mem_init2 = "A9C019559C1CD54E01CAACE0E6AB700CD527DF25598066A93C79AADC03955B80E4AD8FE25523FCCAB60836A91FE35563FCCAB70066AD8FE65533F8DAB30076A91FF36B670E254CFFCD748FE36A4E0396D31E1B54C7F32A99FE65531F8DA930036AB3839B4B1FC6D49C03256CFF9B52600C95B3FE6559803B549F7CD54C7E36A4C00CAADC03B55B8076AA60066AD9FE36A4C019AA4F0E2D68E1E4AB30064AD9FF12A99FE65567FE255B06192D3003356CFF9956C7E36A99FF32AD8FC6D533FE65531F8CAACF9E692CFFC4AB70C3256C7F1B56E3C32AB381C956E006554C00ED56601CB5B3FF36A4C01CB491FC65523FF349670736A4E0392A4C019AADC00CAA98";
defparam ram_block1a120.mem_init1 = "F8ED5B3FE25567039AA98FC6556E00C952701C952600ED54CFF32DA60076AB7003252C7FCDAB63F8DAA67FE6D5B1FC6D5B3FF36AD8FE32A93C1CD259C1E4AA63F8CAA4E0736B6E019B4B383C954C7F9955980335531FC6D533C79A5A70066AB63F192B67DF34B4C0065A59F3CCAB63FC49499FE34AD9FF8D65380192A4E01C95661C32549C0736B4E00ED759F3E4AACE019AAB3C1CDA931F8CA299FF125247FCCAAD87864AD9C0E6D498FC64AD9C0E6D498FC64AD9C0E6D499FE36AB300192A4C0064AB71F8C95B381E4AA678F12AB30033552783C9559801DA4B3007255B1FF32D2C7FF34A58FFC4AA98FE32569C01C956C7FE6D52600335533C7894531FE36";
defparam ram_block1a120.mem_init0 = "AB31F8C956C7F8CA6B3C1E69491FF996D6783895531FE36AA67FF32AA63FE64AD98019A4A61F8C95267FC6D56C7FC6D56C7FCCD56C7FC6D56C7FE65359C0392AB63FC64A930FC64AB63FF1B5498FE3255B3FFCCAAD9FFC695261F0C956CF8F1252CC00E4AACC7E196A48FFE65359C01CD6533FF8DAAD8FFC6D54CE039B55B1FF8DAAD9C0732AA67878D2A4C7F8C956CF03CD29660C19AAB63FF1B552700392AB67FF892A4CFFE36AB6700E6556CF879955270019B56DC3C336A59800E4AA99C079A5499FFE6535B1FF8DAAB63FF992AD9800CCAAD9C038955663F865AA4C7FC65AB6E1F0CD55270039B54B1C0F32D699F0F32D691C039955663FE3255263FF19";

cyclonev_ram_block ram_block1a144(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a144_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a144.clk0_core_clock_enable = "ena0";
defparam ram_block1a144.clk0_input_clock_enable = "ena0";
defparam ram_block1a144.clk0_output_clock_enable = "ena0";
defparam ram_block1a144.data_interleave_offset_in_bits = 1;
defparam ram_block1a144.data_interleave_width_in_bits = 1;
defparam ram_block1a144.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a144.init_file_layout = "port_a";
defparam ram_block1a144.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a144.operation_mode = "rom";
defparam ram_block1a144.port_a_address_clear = "none";
defparam ram_block1a144.port_a_address_width = 13;
defparam ram_block1a144.port_a_data_out_clear = "none";
defparam ram_block1a144.port_a_data_out_clock = "clock0";
defparam ram_block1a144.port_a_data_width = 1;
defparam ram_block1a144.port_a_first_address = 49152;
defparam ram_block1a144.port_a_first_bit_number = 0;
defparam ram_block1a144.port_a_last_address = 57343;
defparam ram_block1a144.port_a_logical_ram_depth = 65536;
defparam ram_block1a144.port_a_logical_ram_width = 24;
defparam ram_block1a144.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a144.ram_block_type = "auto";
defparam ram_block1a144.mem_init3 = "31FF8C95498FF8CD553380712D699E1F32D699E071A55B3801C955661F0EDAB4C7FC64AB4C3F8CD552380736AA6600336A933FF8DAAB63FF1B594CFFF3254B3C0732AA4E00334AD987876D5B3001C95533C3E6D54CE01CDAAD8FFE64A923FFCDAA93801C955B1FF8DAAB3060CD296781E6D5263FC64A963C3CCAA99C0736AB63FF1B55B380E6556C7FE36AB63FF994D670073594CFFE24AD30FC66AA4E00669491E3E6D5261F0C952C7FF36AA67FF9B5498FE3255B1FF8DAA4C7E192A4C7F8DAA938073594CFFC6D56C7FC6D5667FC6D56C7FC6D56C7FCC95263F0CA4B300336A4CFF8CAA99FFCCAAD8FF19552383CD6D33FF1252CF079ACA63FC6D5263F19AA";
defparam ram_block1a144.mem_init2 = "D8FF194523C799559800C956CFFC6D5270072D498FE32AA47FE34A59FFC69699FF1B549C019A4B70033552783C95598019AA91E3CCAA4F039B5263F1DAA4C0064A930019AAD8FF3256CE0736A4C7E3256CE0736A4C7E3256CE0736A4C3C36AA67FC49491FF328A63F192B67079AAB300E6AA4F9F35D6E00E5AD9C072549870CD52700E4A9300394D63FF36A58FF325247F8DAA679F34B4C0065A59F7CDA931F8DAACC01CB4B3C79956C7F1955980335533FC65527839A5B300EDAD9C0E4AA63F8CAA4F07349670792A98FE36AD9FF9B56C7F1B56CFFCCAB63F8DAB67FC6949801DAADC00CB699FE6556E00C952701C952600ED54C7E32AB381CD548FF9B56E3E";
defparam ram_block1a144.mem_init1 = "32AA60076AB30064A9380E4AD9C1CD259FF8954C7F125A70064AD9FF9B5A700CD56E006554C00ED527039AA9878ED5B1FC6D49861DAA47FE692CF3E6AA63F1954CFF9956C7E36A99FF32AD8FC6D533FE6D5980196930C1B548FFCD54CFF32A91FF36A4C019AA4F0E2D68E1E4AB30064AD8FF36ACC00CAADC03B55B8076AA60064AD8FC65567DF255B803354CFF9B52600C95B3FE6D49807256C7F1A5B3839AAD80192B63F1954CFF32A99FC655B0F196D380E4AD8FE25D67FE6548E1CDAD9FF12ADC019AB63F9954CFE36ACC01DAA67F8D558FF12AD820DAA67F89548FE36A4E03B5538076AB3C792ACC033549F7C956601DAACE0E6AA700E55670735530072A";
defparam ram_block1a144.mem_init0 = "B3C79AACE07256C7F12A91FC6D69E1E4AD9FF36B67FE6AA60064A4C0192B61C32CB38792A67FCCA93C39AA982192D380ED56E0396930032AB3EF36B63F8D548FE34B67FE6AB700E5567DE6D6CFF9A4B3FE6D6CF7CD56E01DAA47F8954C00C9498072AB701DAA9C072D26006D533F8DA93C39B498F192D381C95B3FC4AA60064A4E03B559C1CD5278F2548FF89523FE2549FFC95278F3559C1CD56E0396D30066AD820DAA63E32AB1FE6D6CFF895278F3559C0ED54E0396930064A4C019AB70076ADC01DAB70066A4C01929380E5567073549FF9B4B1FCCAB6006596707256C7F32ACC03354CFF32ACC03256C7E34B67FE6AB701C949801B54C7C65523F8D558F";

cyclonev_ram_block ram_block1a168(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a168_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a168.clk0_core_clock_enable = "ena0";
defparam ram_block1a168.clk0_input_clock_enable = "ena0";
defparam ram_block1a168.clk0_output_clock_enable = "ena0";
defparam ram_block1a168.data_interleave_offset_in_bits = 1;
defparam ram_block1a168.data_interleave_width_in_bits = 1;
defparam ram_block1a168.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a168.init_file_layout = "port_a";
defparam ram_block1a168.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a168.operation_mode = "rom";
defparam ram_block1a168.port_a_address_clear = "none";
defparam ram_block1a168.port_a_address_width = 13;
defparam ram_block1a168.port_a_data_out_clear = "none";
defparam ram_block1a168.port_a_data_out_clock = "clock0";
defparam ram_block1a168.port_a_data_width = 1;
defparam ram_block1a168.port_a_first_address = 57344;
defparam ram_block1a168.port_a_first_bit_number = 0;
defparam ram_block1a168.port_a_last_address = 65535;
defparam ram_block1a168.port_a_logical_ram_depth = 65536;
defparam ram_block1a168.port_a_logical_ram_width = 24;
defparam ram_block1a168.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a168.ram_block_type = "auto";
defparam ram_block1a168.mem_init3 = "3C3C3C3C3C3C1E1E0F0F87C1E0F83E0FC1F81F81FC07F007FC00FFFC00001FFFFFFFC00007FF803FC07E07C1F0F0F0E1C78E31CE319CCC66666CC99364924925B4B5AD6A55AA9555555554AAD5A94A5A4B6DB64D9B333399CE31C38787C0FF0007FFC001FC0F87871C6319CCD9936DB69294AD54AAAAB552B5A5A49364CCCC671C70F83F80000001FC1E1C31CC666CDB6DA52954AAAA55294B6DB2666631C787C07FFFFF01F0E18E66664DA4B5AA55556AD696DB327338E1E0FFC01FF83C38C6666C96D6A555556A5A49B33318F0F801FC00F871CE66C925AD55A554A5B6CCCC6387E000007E1C73332692952AA952D24D98C71E07FFFC0F0E73324969555552";
defparam ram_block1a168.mem_init2 = "96C9998E3C07FFC078E33336D2B5555A96D9998E1F00001F0E3333696A555A96933338F03FFE03C63336D295554A5B267387C0000F0E7326D2B555A92C99CF1FC007E1C666DA52AAB5A4998E3C00007863324B5AAA5693633C7F00FE1CE6C96B554A5B6631E00E01E39992D6AAB5A4CCE3C0000F0CCC929555ADB67383FFFE1C666D2AD2ADB6671F0003E399B695556B64E70FE1FE38CDB4AAAA5B66387FFF871992D6AB5A4CC70FFFE1CE4DA5554B6CC70FFFE1C66DAD55293630F001F0CCDB52A56D99C7C01F8E6494AAB49338F801F1CC92955ADB31C1FF838C9A555524CC78000F19B69554B6671FFFF1CCDA5552DB38F803E39B2D554B66707FF0E324B5";
defparam ram_block1a168.mem_init1 = "56926383FE1E66D2AAB6CCE1FFE1CCDA555A4CC7C01F199A555693387FFC31B2D5569B187FFC7336B54A4CC7800F1996A4A9331C001E724A54A4CC7801E33252A52663E01E3934AA96CC700079996AA96CC7C07C724A54A4CE1FFC31B6AAAD99C3FC1CC96AA5B31F83F19B4AAD2638001E649554939E0078CDAD4A4CE3FF87369552CCE07838DB55524E3FFF1C9296A4CE0FC1CC95B52461FFC3325552CC7003C64B55A4C7001E76D55499C3F831B4AA5B387FC3325556CC7C1F19A555B638007992AAB6E7803CCDAAA598F87E725AA5B387F0664AAA4CE060732D55B63800F325556CE3FF0CDAD29338007134AB49C7FF8CDAAAD98FFF8C96A96678078C9554";
defparam ram_block1a168.mem_init0 = "99C003992AADB1F07CCDAAB6E7C1F3B6AADB9F078CD2AD270FF0CCA52998FFC724AA598FFF19B556CC7FF8C96A53380031255499C0073255699E00E3695ACC7FF8CD2A5B1E03C4D6949C7FC324AB4CE003996A9663FF1C95D498FFE336AA4CE00732556DC7FF192AAD9C00312556CC3F866D55B3800734AAD9C081995549C7F866952CC7FE334A9661FC336AA4CF87CC955261FF19B55B30FE19A5693838336AAD8E01C6D55B300066555B3C038DAAB678079B556CE00312D693800725AD23001CDAA931FFC6D296C7FF192A9238073254B31FE336A93380F32D4B3070725549C7E1DB55B3801CD2A59C007255599FFCED6527001CD2B4CF07992ADB87C334AD";

cyclonev_ram_block ram_block1a48(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a48_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a48.clk0_core_clock_enable = "ena0";
defparam ram_block1a48.clk0_input_clock_enable = "ena0";
defparam ram_block1a48.clk0_output_clock_enable = "ena0";
defparam ram_block1a48.data_interleave_offset_in_bits = 1;
defparam ram_block1a48.data_interleave_width_in_bits = 1;
defparam ram_block1a48.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a48.init_file_layout = "port_a";
defparam ram_block1a48.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a48.operation_mode = "rom";
defparam ram_block1a48.port_a_address_clear = "none";
defparam ram_block1a48.port_a_address_width = 13;
defparam ram_block1a48.port_a_data_out_clear = "none";
defparam ram_block1a48.port_a_data_out_clock = "clock0";
defparam ram_block1a48.port_a_data_width = 1;
defparam ram_block1a48.port_a_first_address = 16384;
defparam ram_block1a48.port_a_first_bit_number = 0;
defparam ram_block1a48.port_a_last_address = 24575;
defparam ram_block1a48.port_a_logical_ram_depth = 65536;
defparam ram_block1a48.port_a_logical_ram_width = 24;
defparam ram_block1a48.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a48.ram_block_type = "auto";
defparam ram_block1a48.mem_init3 = "31FF8C95498FF8CD553380712D699E1F32D699E071A55B3801C955661F0EDAB4C7FC64AB4C3F8CD552380736AA6600336A933FF8DAAB63FF1B594CFFF3254B3C0732AA4E00334AD987876D5B3001C95533C3E6D54CE01CDAAD8FFE64A923FFCDAA93801C955B1FF8DAAB3060CD296781E6D5263FC64A963C3CCAA99C0736AB63FF1B55B380E6556C7FE36AB63FF994D670073594CFFE24AD30FC66AA4E00669491E3E6D5261F0C952C7FF36AA67FF9B5498FE3255B1FF8DAA4C7E192A4C7F8DAA938073594CFFC6D56C7FC6D5667FC6D56C7FC6D56C7FCC95263F0CA4B300336A4CFF8CAA99FFCCAAD8FF19552383CD6D33FF1252CF079ACA63FC6D5263F19AA";
defparam ram_block1a48.mem_init2 = "D8FF194523C799559800C956CFFC6D5270072D498FE32AA47FE34A59FFC69699FF1B549C019A4B70033552783C95598019AA91E3CCAA4F039B5263F1DAA4C0064A930019AAD8FF3256CE0736A4C7E3256CE0736A4C7E3256CE0736A4C3C36AA67FC49491FF328A63F192B67079AAB300E6AA4F9F35D6E00E5AD9C072549870CD52700E4A9300394D63FF36A58FF325247F8DAA679F34B4C0065A59F7CDA931F8DAACC01CB4B3C79956C7F1955980335533FC65527839A5B300EDAD9C0E4AA63F8CAA4F07349670792A98FE36AD9FF9B56C7F1B56CFFCCAB63F8DAB67FC6949801DAADC00CB699FE6556E00C952701C952600ED54C7E32AB381CD548FF9B56E3E";
defparam ram_block1a48.mem_init1 = "32AA60076AB30064A9380E4AD9C1CD259FF8954C7F125A70064AD9FF9B5A700CD56E006554C00ED527039AA9878ED5B1FC6D49861DAA47FE692CF3E6AA63F1954CFF9956C7E36A99FF32AD8FC6D533FE6D5980196930C1B548FFCD54CFF32A91FF36A4C019AA4F0E2D68E1E4AB30064AD8FF36ACC00CAADC03B55B8076AA60064AD8FC65567DF255B803354CFF9B52600C95B3FE6D49807256C7F1A5B3839AAD80192B63F1954CFF32A99FC655B0F196D380E4AD8FE25D67FE6548E1CDAD9FF12ADC019AB63F9954CFE36ACC01DAA67F8D558FF12AD820DAA67F89548FE36A4E03B5538076AB3C792ACC033549F7C956601DAACE0E6AA700E55670735530072A";
defparam ram_block1a48.mem_init0 = "B3C79AACE07256C7F12A91FC6D69E1E4AD9FF36B67FE6AA60064A4C0192B61C32CB38792A67FCCA93C39AA982192D380ED56E0396930032AB3EF36B63F8D548FE34B67FE6AB700E5567DE6D6CFF9A4B3FE6D6CF7CD56E01DAA47F8954C00C9498072AB701DAA9C072D26006D533F8DA93C39B498F192D381C95B3FC4AA60064A4E03B559C1CD5278F2548FF89523FE2549FFC95278F3559C1CD56E0396D30066AD820DAA63E32AB1FE6D6CFF895278F3559C0ED54E0396930064A4C019AB70076ADC01DAB70066A4C01929380E5567073549FF9B4B1FCCAB6006596707256C7F32ACC03354CFF32ACC03256C7E34B67FE6AB701C949801B54C7C65523F8D558F";

cyclonev_ram_block ram_block1a72(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a72_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a72.clk0_core_clock_enable = "ena0";
defparam ram_block1a72.clk0_input_clock_enable = "ena0";
defparam ram_block1a72.clk0_output_clock_enable = "ena0";
defparam ram_block1a72.data_interleave_offset_in_bits = 1;
defparam ram_block1a72.data_interleave_width_in_bits = 1;
defparam ram_block1a72.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a72.init_file_layout = "port_a";
defparam ram_block1a72.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a72.operation_mode = "rom";
defparam ram_block1a72.port_a_address_clear = "none";
defparam ram_block1a72.port_a_address_width = 13;
defparam ram_block1a72.port_a_data_out_clear = "none";
defparam ram_block1a72.port_a_data_out_clock = "clock0";
defparam ram_block1a72.port_a_data_width = 1;
defparam ram_block1a72.port_a_first_address = 24576;
defparam ram_block1a72.port_a_first_bit_number = 0;
defparam ram_block1a72.port_a_last_address = 32767;
defparam ram_block1a72.port_a_logical_ram_depth = 65536;
defparam ram_block1a72.port_a_logical_ram_width = 24;
defparam ram_block1a72.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a72.ram_block_type = "auto";
defparam ram_block1a72.mem_init3 = "3C3C3C3C3C3C1E1E0F0F87C1E0F83E0FC1F81F81FC07F007FC00FFFC00001FFFFFFFC00007FF803FC07E07C1F0F0F0E1C78E31CE319CCC66666CC99364924925B4B5AD6A55AA9555555554AAD5A94A5A4B6DB64D9B333399CE31C38787C0FF0007FFC001FC0F87871C6319CCD9936DB69294AD54AAAAB552B5A5A49364CCCC671C70F83F80000001FC1E1C31CC666CDB6DA52954AAAA55294B6DB2666631C787C07FFFFF01F0E18E66664DA4B5AA55556AD696DB327338E1E0FFC01FF83C38C6666C96D6A555556A5A49B33318F0F801FC00F871CE66C925AD55A554A5B6CCCC6387E000007E1C73332692952AA952D24D98C71E07FFFC0F0E73324969555552";
defparam ram_block1a72.mem_init2 = "96C9998E3C07FFC078E33336D2B5555A96D9998E1F00001F0E3333696A555A96933338F03FFE03C63336D295554A5B267387C0000F0E7326D2B555A92C99CF1FC007E1C666DA52AAB5A4998E3C00007863324B5AAA5693633C7F00FE1CE6C96B554A5B6631E00E01E39992D6AAB5A4CCE3C0000F0CCC929555ADB67383FFFE1C666D2AD2ADB6671F0003E399B695556B64E70FE1FE38CDB4AAAA5B66387FFF871992D6AB5A4CC70FFFE1CE4DA5554B6CC70FFFE1C66DAD55293630F001F0CCDB52A56D99C7C01F8E6494AAB49338F801F1CC92955ADB31C1FF838C9A555524CC78000F19B69554B6671FFFF1CCDA5552DB38F803E39B2D554B66707FF0E324B5";
defparam ram_block1a72.mem_init1 = "56926383FE1E66D2AAB6CCE1FFE1CCDA555A4CC7C01F199A555693387FFC31B2D5569B187FFC7336B54A4CC7800F1996A4A9331C001E724A54A4CC7801E33252A52663E01E3934AA96CC700079996AA96CC7C07C724A54A4CE1FFC31B6AAAD99C3FC1CC96AA5B31F83F19B4AAD2638001E649554939E0078CDAD4A4CE3FF87369552CCE07838DB55524E3FFF1C9296A4CE0FC1CC95B52461FFC3325552CC7003C64B55A4C7001E76D55499C3F831B4AA5B387FC3325556CC7C1F19A555B638007992AAB6E7803CCDAAA598F87E725AA5B387F0664AAA4CE060732D55B63800F325556CE3FF0CDAD29338007134AB49C7FF8CDAAAD98FFF8C96A96678078C9554";
defparam ram_block1a72.mem_init0 = "99C003992AADB1F07CCDAAB6E7C1F3B6AADB9F078CD2AD270FF0CCA52998FFC724AA598FFF19B556CC7FF8C96A53380031255499C0073255699E00E3695ACC7FF8CD2A5B1E03C4D6949C7FC324AB4CE003996A9663FF1C95D498FFE336AA4CE00732556DC7FF192AAD9C00312556CC3F866D55B3800734AAD9C081995549C7F866952CC7FE334A9661FC336AA4CF87CC955261FF19B55B30FE19A5693838336AAD8E01C6D55B300066555B3C038DAAB678079B556CE00312D693800725AD23001CDAA931FFC6D296C7FF192A9238073254B31FE336A93380F32D4B3070725549C7E1DB55B3801CD2A59C007255599FFCED6527001CD2B4CF07992ADB87C334AD";

cyclonev_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 8191;
defparam ram_block1a0.port_a_logical_ram_depth = 65536;
defparam ram_block1a0.port_a_logical_ram_width = 24;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init3 = "6A5987C3B6A933C1E65A967001C94D6E7FF335549C00734A9670039B55B70FC725549C1C19A5699E03992AD98FF19A5499C03892A931FFC6D296C7FF192AB67001896B49C00392D691800E6D55B3C03CDAAB638079B554CC0019B556C700E36AAD9838392D4B30FE19B55B31FF0C955267C3E64AAD987F0CD2A598FFC66952CC3FC7255533020736AA59C0039B556CC3F866D5491800736AA931FFC76D5499C00E64AAD98FFE32575271FF8CD2AD33800E65AA4987FC7252D64780F1B4A9663FFC66B52D8E00F32D5499C00732554918003994AD263FFC66D55B31FFE334AA49C7FE33294A661FE1C96A9663C1F3B6AADB9F07CEDAAB667C1F1B6AA933800732";
defparam ram_block1a0.mem_init2 = "555263C03CCD2AD263FFE336AAB663FFC725AA591C00399296B661FF8E6D55499E0038DB55699C0C0E64AAA4CC1FC39B4AB49CFC3E334AAB667803CEDAAA933C0038DB554B31F07C66D5549987FC39B4AA5B183F87325556DCF001C64B55A4C7801C6695549987FF0C495B526707E0E64AD29271FFF8E49555B6383C0E669552D9C3FF8E64A56B663C00F39255524CF00038C96AA5B31F83F19B4AAD26707F87336AAADB187FF0E64A54A49C7C07C66D2AAD333C001C66D2AA5938F00F8CC94A94998F003C664A54A49CF00071992A4AD331E003C664A55AD99C7FFC31B2D5569B187FFC3992D554B331F007C664B554B6670FFF0E66DAAA96CCF0FF838C92D5";
defparam ram_block1a0.mem_init1 = "5A498E1FFC1CCDA55569B38F803E39B69554B6671FFFF1CCDA5552DB31E0003C66495554B26383FF0719B6B55292671F003E39925AAA524CE3F007C7336D4A95B6661F001E18D929556B6CC70FFFE1C66DA5554B64E70FFFE1C664B5AAD69331C3FFFC38CDB4AAAA5B6638FF0FE1CE4DAD5552DB338F8001F1CCDB6A96A96CCC70FFFF839CDB6B5552926661E000078E664B5AAAD693338F00E00F18CDB4A555AD26CE70FE01FC798D92D4AAB5A4998C3C000078E3324B5AAA94B6CCC70FC007F1E732692B555A96C99CE1E00007C39CC9B4A5555296D998C780FFF81E399992D2B554AD2D9998E1F00001F0E33336D2B5555A96D9998E3C07FFC078E33326D2";
defparam ram_block1a0.mem_init0 = "9555552D24999CE1E07FFFC0F1C6336496952AA95292C9999C70FC00000FC38C6666DB4A554B556B4926CCE71C3E007F003E1E31999B24B4AD55554AD6D26CCCC638783FF007FE0F0E399C99B6D2D6AD5554AB5A4B64CCCCE30E1F01FFFFFC07C3C718CCCC9B6DA52954AAAA55294B6DB66CCC671870F07F00000003F83E1C71CC66664D924B4B5A955AAAAA556A5292DB6D933667318C71C3C3E07F0007FFC001FE07C3C38718E7339999B364DB6DA4B4A52B56AA5555555552AB54AD6B5A5B4924924D93266CCCCC667318E718E3C70E1E1E1F07C0FC07F803FFC00007FFFFFFF000007FFE007FC01FC07F03F03F07E0F83E0F07C3E1E0F0F0787878787878";

cyclonev_ram_block ram_block1a24(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.clk0_output_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "rom";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "clock0";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 8192;
defparam ram_block1a24.port_a_first_bit_number = 0;
defparam ram_block1a24.port_a_last_address = 16383;
defparam ram_block1a24.port_a_logical_ram_depth = 65536;
defparam ram_block1a24.port_a_logical_ram_width = 24;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init3 = "E35563F8954C7C655B003252701DAACFFCDA58FC6D498066A99FE65598066A99FC6D49C1CD34C00DAA67F1A5B3FF2559C1CD54E0392930064ACC01DAB70076ADC01DAB30064A4C0192D380E556E073559E3C9523FE6D6CFF1AA98F8CAB60836ACC0196D380ED567073559E3C9527FF2548FF89523FE2549E3C956707355B80E4A4C00CAA47F9B5270396931E325B38792B63F9956C00C969C072AB701DAA9C0325260065523FC4AB700ED567DE6D6CFF9A4B3FE6D6CF7CD54E01DAACFFCDA58FE25563F8DAD9EF9AA980192D380ED56E0396930832AB38792A67FCCA93C39A69870DA930064A4C00CAACFFCDAD9FF36A4F0F2D6C7F12A91FC6D49C0E6AB3C79A";
defparam ram_block1a24.mem_init2 = "A9C019559C1CD54E01CAACE0E6AB700CD527DF25598066A93C79AADC03955B80E4AD8FE25523FCCAB60836A91FE35563FCCAB70066AD8FE65533F8DAB30076A91FF36B670E254CFFCD748FE36A4E0396D31E1B54C7F32A99FE65531F8DA930036AB3839B4B1FC6D49C03256CFF9B52600C95B3FE6559803B549F7CD54C7E36A4C00CAADC03B55B8076AA60066AD9FE36A4C019AA4F0E2D68E1E4AB30064AD9FF12A99FE65567FE255B06192D3003356CFF9956C7E36A99FF32AD8FC6D533FE65531F8CAACF9E692CFFC4AB70C3256C7F1B56E3C32AB381C956E006554C00ED56601CB5B3FF36A4C01CB491FC65523FF349670736A4E0392A4C019AADC00CAA98";
defparam ram_block1a24.mem_init1 = "F8ED5B3FE25567039AA98FC6556E00C952701C952600ED54CFF32DA60076AB7003252C7FCDAB63F8DAA67FE6D5B1FC6D5B3FF36AD8FE32A93C1CD259C1E4AA63F8CAA4E0736B6E019B4B383C954C7F9955980335531FC6D533C79A5A70066AB63F192B67DF34B4C0065A59F3CCAB63FC49499FE34AD9FF8D65380192A4E01C95661C32549C0736B4E00ED759F3E4AACE019AAB3C1CDA931F8CA299FF125247FCCAAD87864AD9C0E6D498FC64AD9C0E6D498FC64AD9C0E6D499FE36AB300192A4C0064AB71F8C95B381E4AA678F12AB30033552783C9559801DA4B3007255B1FF32D2C7FF34A58FFC4AA98FE32569C01C956C7FE6D52600335533C7894531FE36";
defparam ram_block1a24.mem_init0 = "AB31F8C956C7F8CA6B3C1E69491FF996D6783895531FE36AA67FF32AA63FE64AD98019A4A61F8C95267FC6D56C7FC6D56C7FCCD56C7FC6D56C7FE65359C0392AB63FC64A930FC64AB63FF1B5498FE3255B3FFCCAAD9FFC695261F0C956CF8F1252CC00E4AACC7E196A48FFE65359C01CD6533FF8DAAD8FFC6D54CE039B55B1FF8DAAD9C0732AA67878D2A4C7F8C956CF03CD29660C19AAB63FF1B552700392AB67FF892A4CFFE36AB6700E6556CF879955270019B56DC3C336A59800E4AA99C079A5499FFE6535B1FF8DAAB63FF992AD9800CCAAD9C038955663F865AA4C7FC65AB6E1F0CD55270039B54B1C0F32D699F0F32D691C039955663FE3255263FF19";

cyclonev_ram_block ram_block1a97(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a97_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a97.clk0_core_clock_enable = "ena0";
defparam ram_block1a97.clk0_input_clock_enable = "ena0";
defparam ram_block1a97.clk0_output_clock_enable = "ena0";
defparam ram_block1a97.data_interleave_offset_in_bits = 1;
defparam ram_block1a97.data_interleave_width_in_bits = 1;
defparam ram_block1a97.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a97.init_file_layout = "port_a";
defparam ram_block1a97.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a97.operation_mode = "rom";
defparam ram_block1a97.port_a_address_clear = "none";
defparam ram_block1a97.port_a_address_width = 13;
defparam ram_block1a97.port_a_data_out_clear = "none";
defparam ram_block1a97.port_a_data_out_clock = "clock0";
defparam ram_block1a97.port_a_data_width = 1;
defparam ram_block1a97.port_a_first_address = 32768;
defparam ram_block1a97.port_a_first_bit_number = 1;
defparam ram_block1a97.port_a_last_address = 40959;
defparam ram_block1a97.port_a_logical_ram_depth = 65536;
defparam ram_block1a97.port_a_logical_ram_width = 24;
defparam ram_block1a97.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a97.ram_block_type = "auto";
defparam ram_block1a97.mem_init3 = "1934AD6ADB31C3FFE1C64D2AAA926E707FF0F3324AAAA593187FFF87336D5A95B6671FE3F86324B5552DB31E0FF079CDB4AAAD24CE3E003E31B252AA524CC7800078E6DB55552498E1FFFE1CCC96AAA96CCC7C00078CCDA55552D998F8001F199B4A92ADB673C0FE078CC96B55A9266387FFE1C664B52A569B39E0FFC1E7365A956A4999C3FDFF0E66CB55552D998F03F81E3324B5555A4CCE3E003F1CCDB4AAAB49331E0FFE0E3136D4AAD69B31C3FFFE1C66DB52A95B64E787FFF0739B2D6AA94B2631F0000F1CCDB4AAAA5B6671E000078C64929556B4999C3E001F0C66DB52AB5A4D8C781FE038E64D29555ADB331C1FFFC1C666D2D555ADB331C3FFFF0E";
defparam ram_block1a97.mem_init2 = "3336D6AAA969B31C7C001F0E666D29556A49339E1FFFF8718D92D4AAD4B66671E00007C73324B55954B6CCC70FE03F8739924A5554A593338780003E3999B6955552926673C1FFFC1E33324B52A952D9339C1FC07F0E33324A55556B6D99C707FFFC1E73324B52AA56926C6387F81FE1C636492B5552B6D999C7C03C01E18CC9B4A9552B49367387C0000F8E3336DA555552924CC63C1FFFF078C66492D52AD5A5B3331C1F800FE1C6326DB52AAA94B64CCE3C3FFFFC1E31993495AAAAD6926CE71E0FFFFC1E39CD924A55555AD24C8CE3C1FFFFC1E39CC9B4B52AA95ADB66671C1F8003F871CCCD9694AAAA94B6D998C787F000FE1E3999B25A55AAD5292499";
defparam ram_block1a97.mem_init1 = "9C71F01FFC03C39CCCDB695AAAAB52DB266738781FFFF03C39CCC9B694AAAAA94B6D9998C383FC00FF078E7336492D4AAAAB52DB6CCC638F03FFFFC0F0E339B36D2D4AAAAB52924D998C70F80FFFE03E1C633326D252A5554A94B6D93318E3C1FC0003F83C73999936D295AAAAB56B693666631C3C0FFFFFF03C38E67264DA5AD5AAAAD5296DB266631C787E0000007E1E38C6664DB696A555B555AD6926C999CE38F07F000003F87C71CC666C924B5A95555552B5A4926CCCE738F0F80FFFFFF01F0E18E733364DA4B5AB5555556AD692D936666318E1E0F800FFF801F87871CE7332649B4B4A54AAAAAAA54A5A5B64D9999CE71E1E0FC007FFC007E0F0E1CE";
defparam ram_block1a97.mem_init0 = "73333364924B4A54AAD5556AA56B5A4924D9B3319CE30E1E1F80FFFFFFFFC07C1E1E38C633393326DB6DA5AD4A95552A5554AB5AD2D24926C999998CE71C70F0F83F803FFFFFFE00FE0783878E31CE63333266C926D25A5A56A54AAB555556AA956A529696D249364D99333399CE738E3870F0781F80FF800000000007FE03F03C1E1E3C71C738C6733999993326C9B64924B692D294A52B56A9552AAAAD556AAAAB556A952A52B5A52D2D25B6924936D9364D9B3366666666633398CE739C638E38E38E1C3870F0F0787C1F07E0FC07F01FE01FF800FFF80003FFFFFFF80000000FFFFFFFFE00003FFFC000FFF000FFE007FE00FFC01FE00FF007F807F807F8";

cyclonev_ram_block ram_block1a121(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a121_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a121.clk0_core_clock_enable = "ena0";
defparam ram_block1a121.clk0_input_clock_enable = "ena0";
defparam ram_block1a121.clk0_output_clock_enable = "ena0";
defparam ram_block1a121.data_interleave_offset_in_bits = 1;
defparam ram_block1a121.data_interleave_width_in_bits = 1;
defparam ram_block1a121.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a121.init_file_layout = "port_a";
defparam ram_block1a121.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a121.operation_mode = "rom";
defparam ram_block1a121.port_a_address_clear = "none";
defparam ram_block1a121.port_a_address_width = 13;
defparam ram_block1a121.port_a_data_out_clear = "none";
defparam ram_block1a121.port_a_data_out_clock = "clock0";
defparam ram_block1a121.port_a_data_width = 1;
defparam ram_block1a121.port_a_first_address = 40960;
defparam ram_block1a121.port_a_first_bit_number = 1;
defparam ram_block1a121.port_a_last_address = 49151;
defparam ram_block1a121.port_a_logical_ram_depth = 65536;
defparam ram_block1a121.port_a_logical_ram_width = 24;
defparam ram_block1a121.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a121.ram_block_type = "auto";
defparam ram_block1a121.mem_init3 = "1F332952D98F83E336AAA49C7FFC665AA96C60FC1CDB554B31E01E334AAB4CE1FC1CDB5569B8FFFC66D2A5363C00E334AA966700071B6AAB6CF0003992AAA4CE0003996AAB6C700071B6AAB667000F334AA9263C01E325AA5331F07C66D5D5B30FFF8E495549987FF0CCB556D9C7FF1CDA552D9C3FE1CDB556D987FF0CC9554938FFFC66D2AD26380071B6B4A49C3FF8E6D6AD26700038DB555B33800399B555B638001CC96A96CC7FFE332D54B670FF8626954B670FFC3325556CCF003C6CA54B667C07C64B552CCE00071B6AAB66700071B6A2A4CC3FF8E6D2A96CE3FF8624ADA931C001C6DAAA9330FFC39B4AA5B38FFF1CDAD5A4CE1FC1CDB554B33C0079";
defparam ram_block1a121.mem_init2 = "9B5552661FFC3325556CCF001E66D55699C7FF1CCB554B31C00799B5552663FFE39B5AB499C3FC3992A2A4CE1FE0CCD6A96CC7FFE19B5AB499C3F83996AAA4CE1FF0E6D2AB498F003CEDA54A4C700071B6B4AD98F80F19B4AB499C1F839B6AAA4CC3FF8726B56B671FFF1CDA552D9C7FFC736954B661FFF8CDB556998F81F1925556CCE0007336AAA4CC7FFE19B4AB5B38FFF866DAAB498F001C669554931E00F19B4AB49987FE1CC953524E3FFF0CDA552D98F81F19B4AA5B31F03E336954B663E07C665AAB4DCF003C66D595B6707F07325695B33C0038CDAAAB6670001CCD2AA9263C00F1925556D8E1FC1CC96AA59187FF0E6DAAADB38FFF8664AAA9331F";
defparam ram_block1a121.mem_init1 = "07E336954B667800799B5A94998FFFC736D556D9C7FFE3325AA5B638000E66D555B6307FC399295293387FE1CC94A9499C3FF0E64A54A4CE3FFC3134AAB6CC7C07C66DAAA5B38FFF87269556D98F8078CCB555A663E03E3369552C9C7FFE199295ADB387FF0C6DAAAB6C61FFC39929569271E01F39B4AAD6463FFF8E6DAAA926781C0E324AAA5B38FFFE3134AAB6CCF00079996AA96CE3E07C664B55A49C7803C664AD2B6CE1FFE1CDB5A94931E001E324A56B6CE1FFE1CDB4AB5B33C0007192555493381F838C96AAB6CC7800F1996AAA599C7FFC7334AAA9373C000E336B55A49CF800F3935AA96CCE0FE0E324AAA926707FE1CC92AAA599C3FF87336B54A4";
defparam ram_block1a121.mem_init0 = "CC3E07C73252AD6C8C3FFE18DB4AAD24E780078CC94AB5B3387FF0E66D6AB4931E00079D92B52926387FC1CCDAD56B66707FC3CCDAD56B66707FE1CECB55524CC7C03E39B6A56B6CC7C00F8CDB5AB5B663C003C664B556B26381F038CDA555A49CF0001C665AD4ADB38F001E3134AAA96463C007C664A556B6670FFF87336B5529331E000F1992D5529B38F807C7325AAA964E780C079992955AD99C7FFF8E66D2AAD24C70FFE0E66D2AAB4998F00078CC92AAAD2671FC3F0E6CB55549331E00079CDB4AAB49B9C1FF8399929552DB31E0003C664B5552D9987C07E399252A949338FE0FC3336D5552D98C1FFF0E324B555A498E1FFF87332D6AB5B66383FF07";

cyclonev_ram_block ram_block1a145(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a145_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a145.clk0_core_clock_enable = "ena0";
defparam ram_block1a145.clk0_input_clock_enable = "ena0";
defparam ram_block1a145.clk0_output_clock_enable = "ena0";
defparam ram_block1a145.data_interleave_offset_in_bits = 1;
defparam ram_block1a145.data_interleave_width_in_bits = 1;
defparam ram_block1a145.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a145.init_file_layout = "port_a";
defparam ram_block1a145.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a145.operation_mode = "rom";
defparam ram_block1a145.port_a_address_clear = "none";
defparam ram_block1a145.port_a_address_width = 13;
defparam ram_block1a145.port_a_data_out_clear = "none";
defparam ram_block1a145.port_a_data_out_clock = "clock0";
defparam ram_block1a145.port_a_data_width = 1;
defparam ram_block1a145.port_a_first_address = 49152;
defparam ram_block1a145.port_a_first_bit_number = 1;
defparam ram_block1a145.port_a_last_address = 57343;
defparam ram_block1a145.port_a_logical_ram_depth = 65536;
defparam ram_block1a145.port_a_logical_ram_width = 24;
defparam ram_block1a145.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a145.ram_block_type = "auto";
defparam ram_block1a145.mem_init3 = "C1FF838CDB5AAD6999C3FFF0E324B555A498E1FFF0633695556D9987E0FE399252A949338FC07C33369555A4CC78000F19B69552933383FF073B25AAA5B673C000F19925555A6CE1F87F1CC96AAA92663C001E3325AAA96CCE0FFE1C6496AA96CCE3FFFC7336B5529333C0603CE4D2AAB499C7C03E39B295569331E000F1992955AD99C3FFE1CCDAD54A4CC7C0078C4D2AAA5918F001E39B6A56B4CC70001E724B554B66381F038C9AD55A4CC780078CDB5AB5B663E007C66DAD4ADB38F807C6649555A6E70FFC1CCDAD56B66787FC1CCDAD56B66707FC38C9295A9373C000F1925AAD6CCE1FFC399B5AA52663C003CE496AA5B630FFF8626D6A9499C7C0F866";
defparam ram_block1a145.mem_init2 = "4A55AD99C3FF87334AAA92670FFC1CC92AAA498E0FE0E66D2AB5939E003E724B55AD98E00079D92AAA599C7FFC7334AAAD331E003C66DAAAD26383F039925554931C000799B5AA5B670FFF0E6DAD4A498F000F19252B5B670FFF0E6DA96A4CC7803C724B55A4CC7C0F8E6D2AAD333C001E66DAAA5918FFFE39B4AAA498E0703CC92AAB6CE3FFF8C4D6AA5B39F00F1C92D5293387FF0C6DAAAB6C61FFC39B6B529330FFFC7269552D98F80F8CCB555A663C03E336D552C9C3FFE39B4AAB6CC7C07C66DAAA59187FF8E64A54A4CE1FF873252A52670FFC399295293387FC18DB5556CCE00038DB4AB4998FFFC736D556D9C7FFE33252B5B33C003CCDA552D98FC1";
defparam ram_block1a145.mem_init1 = "F1992AAA4CC3FFE39B6AAB6CE1FFC3134AAD26707F0E36D554931E0078C92AA96670001CCDAAAB663800799B52D499C1FC1CDB5356CC7801E765AAB4CC7C0F8CDA552D98F81F19B4AA5B31F03E336954B661FFF8E495952670FFC3325AA5B31E00F1925552CC7001E325AAB6CC3FFE39B5AA5B30FFFC664AAAD99C000E66D554931F03E332D55B663FFF0CDA552D9C7FFC736954B671FFF1CDAD5AC9C3FF8664AAADB383F07325AA5B31E03E336A5ADB1C001C64A54B6E7801E325AA96CE1FF0E64AAAD3383F87325AB5B30FFFC66D2AD6660FF0E64A8A93387F87325AB5B38FFF8CC9555B33C00719A555A671FFC732D556CCF001E66D5549987FF0CC9555B3";
defparam ram_block1a145.mem_init0 = "3C00799A555B6707F0E64B56B671FFE39B4AA5B387FE1992AAB6C70007192B6A48C3FF8E6D2A96CE3FF8664A8ADB1C001CCDAAADB1C000E66955A4C7C07CCDA54A6C7801E66D5549987FE1CDA552C8C3FE1CDA556998FFFC66D2AD26700038DB555B33800399B555B638001CC96AD6CE3FF8724A5ADB1C0038C96A96CC7FFE3925552661FFC336D55B670FF8736954B671FFC736D55A661FFC33255524E3FFE19B5756CC7C1F1994AB498F0078C92AA599E001CCDAAADB1C001C6DAAAD338000E64AAA9338001E6DAAADB1C001CCD2AA598E0078D94A96CC7FFE3B2D55B6707F0E65AAA598F00F19A555B6707E0C6D2AB4CC7FFC724AAAD98F83E336952999F0";

cyclonev_ram_block ram_block1a169(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a169_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a169.clk0_core_clock_enable = "ena0";
defparam ram_block1a169.clk0_input_clock_enable = "ena0";
defparam ram_block1a169.clk0_output_clock_enable = "ena0";
defparam ram_block1a169.data_interleave_offset_in_bits = 1;
defparam ram_block1a169.data_interleave_width_in_bits = 1;
defparam ram_block1a169.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a169.init_file_layout = "port_a";
defparam ram_block1a169.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a169.operation_mode = "rom";
defparam ram_block1a169.port_a_address_clear = "none";
defparam ram_block1a169.port_a_address_width = 13;
defparam ram_block1a169.port_a_data_out_clear = "none";
defparam ram_block1a169.port_a_data_out_clock = "clock0";
defparam ram_block1a169.port_a_data_width = 1;
defparam ram_block1a169.port_a_first_address = 57344;
defparam ram_block1a169.port_a_first_bit_number = 1;
defparam ram_block1a169.port_a_last_address = 65535;
defparam ram_block1a169.port_a_logical_ram_depth = 65536;
defparam ram_block1a169.port_a_logical_ram_width = 24;
defparam ram_block1a169.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a169.ram_block_type = "auto";
defparam ram_block1a169.mem_init3 = "3FC03FC03FC01FE00FF007FE00FFC00FFE001FFE0007FFF80000FFFFFFFFE00000003FFFFFFF80003FFE003FF00FF01FC07E0FC1F07C3C1E1E1C3870E38E38E38C739CE633998CCCCCCCCD99B364D936D92492DB4969694B5A94A952AD55AAAAAD556AAAA9552AD5A94A529692DA4924DB26C9993333399CC639C71C78F0F0781F80FFC00000000003FE03F03C1E1C38E39CE73399993364D92496D2D294AD52AAD55555AAA54AD4B4B496C926CC99998CE718E3C383C0FE00FFFFFFF803F83E1E1C71CE63333326C9249696B5AA5554A95552A56B4B6DB6C9993998C638F0F07C07FFFFFFFE03F0F0E18E73199B364924B5AD4AAD5556AA54A5A4924D99999C";
defparam ram_block1a169.mem_init2 = "E70E1E0FC007FFC007E0F0F1CE7333364DB4B4A54AAAAAAA54A5A5B24C999CE71C3C3F003FFE003E0F0E318CCCD93692D6AD555555AB5A4B64D999CE30E1F01FFFFFE03E1E39CE666C924B5A95555552B5A4926CCC671C7C3F800001FC1E38E73326C92D6B555B554AD2DB64CCC638F0FC000000FC3C718CCC9B6D2956AAAB56B4B64C9CCE38781FFFFFE078718CCCD92DAD5AAAAB5296D933339C783F80007F078E319936DA52A5554A9496C9998C70F80FFFE03E1C6333649295AAAAA5696D9B398E1E07FFFF81E38C666DB695AAAAA56924D99CE3C1FE007F838633336DA52AAAAA52DB266738781FFFF03C39CCC9B695AAAAB52DB6667387807FF01F1C73";
defparam ram_block1a169.mem_init1 = "32492956AB54B49B3338F0FE001FC3C63336DA52AAAA52D366671C3F8003F071CCCDB6B52AA95A5B26738F07FFFF078E626496B55554A4936738F07FFFE0F1CE6C92D6AAAB52593318F07FFFF878E664DA52AAA95B6C98C70FE003F071999B4B56A956924CC63C1FFFF078C66492955554B6D998E3E00007C39CD925A9552A5B26630F007807C73336DA9555A924D8C70FF03FC38C6C92D4AA95A4999CF07FFFC1C7336DAD5554A49998E1FC07F0739936952A95A49998F07FFF079CCC92955552DB3338F80003C399934A5554A49339C3F80FE1C666DA55355A4999C7C0000F1CCCDA56AA5693631C3FFFF0F39924AD55296CCCE1F0007C719B2D2AAAD6D998";
defparam ram_block1a169.mem_init0 = "E1FFFF87199B6B555696CCC707FFF07199B6B5552964CE380FF03C6364B5AA95B6CC61F000F873325AD552924C63C0000F1CCDB4AAAA5B6671E0001F18C9A52AAD69B39C1FFFC3CE4DB52A95B6CC70FFFF8719B2D6AA56D918E0FFE0F19925AAAA5B6671F800F8E664B5555A4998F03F81E333695555A6CCE1FF7F873324AD52B4D9CF07FE0F39B2D4A95A4CC70FFFC38CC92B55AD2663C0FE079CDB6A92A5B331F0003E333695554B6663C0007C666D2AAAD26670FFFF0E32495555B6CE3C0003C66494AA949B18F800F8E6496AAA5B673C1FE0F19B69555A498C3F8FF1CCDB52B56D99C3FFFC31934AAAA4999E1FFC1CEC92AAA964C70FFF8719B6AD6A5931";

cyclonev_ram_block ram_block1a49(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a49_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a49.clk0_core_clock_enable = "ena0";
defparam ram_block1a49.clk0_input_clock_enable = "ena0";
defparam ram_block1a49.clk0_output_clock_enable = "ena0";
defparam ram_block1a49.data_interleave_offset_in_bits = 1;
defparam ram_block1a49.data_interleave_width_in_bits = 1;
defparam ram_block1a49.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a49.init_file_layout = "port_a";
defparam ram_block1a49.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a49.operation_mode = "rom";
defparam ram_block1a49.port_a_address_clear = "none";
defparam ram_block1a49.port_a_address_width = 13;
defparam ram_block1a49.port_a_data_out_clear = "none";
defparam ram_block1a49.port_a_data_out_clock = "clock0";
defparam ram_block1a49.port_a_data_width = 1;
defparam ram_block1a49.port_a_first_address = 16384;
defparam ram_block1a49.port_a_first_bit_number = 1;
defparam ram_block1a49.port_a_last_address = 24575;
defparam ram_block1a49.port_a_logical_ram_depth = 65536;
defparam ram_block1a49.port_a_logical_ram_width = 24;
defparam ram_block1a49.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a49.ram_block_type = "auto";
defparam ram_block1a49.mem_init3 = "F0000F1992D555A4CCF07F81CE4D2B4A964E781F81C66DAD54A4CCE1FFF0E32695552D98C3FFF0E664AD5292661E003C7325AAAA4998E0001C626955569338FC07C3336B556926387FF871925AAB5B330FC3F8E6694AB5B663800078CDB5555B66707FE0E66DAAAA4998F000F1CDB52B524CE1FFF87324A96A59987C07C7324AAAB6CC707F0799B6AAA92671FFFE189B5AAD6C8C3FFFC7365AAAD2663E0078E6DAB6ADB31E000F19B6AAA92661FFFE3992D5569338FFFF1CC96AAB499C3FFF1CCDAD529373C000719B6AAADB31E000719B6AAADB31C000F19B4AAA5938F003C7369555A6678000F336D554B331F83F189A5554931C0F81CECB55524CE1FFE1CC";
defparam ram_block1a49.mem_init2 = "92AAB4DCE0381E66D2AA5B31C000719B5AAD64C78003CCC95556D9C7FFF8E4D2AAB6CC7C01E3925AA96CCE07C0E66D2AB4998FE3F0CC95A94931E001E3369552D98F001E336D556931C1F838C96AA96CE3E07C7369556931C1F838C96AA92661FFF8E6DAAA96461FFE1CDB5AD4998F00F8CC95356CCE1FF0636D6AD6CC7800F19B5AA52670FFC189B5556D9C7FFC39B6AAA499E06038D96AAD3638080E325AAA499C3FE0C6DA92B4CE3FFE1992D569330FFF8664AD6B6C70FF0E36D6A52661FFF0CC95AD6D8E0F81CCD2AA92638001C649554931C000F324AAA498E0007192D54B663C00F3B2D552CCE1FF0E64A54A4CE1FF0E669556998F81F1992AAB6CE1FF";
defparam ram_block1a49.mem_init1 = "C3334AAD2670FF873252A526383E0E36D555B33C001C6CA552D9C7FFE3935AA5B31E0079996AA5B31F03E332D55A4C70007192D54B663FFF8E495952661FFE1996AAB4CE3FFC732D55699C7FF8E65AAADB387FE18DA5549338000E669556998FFFC736954B663F0FCE4D4B52670FF8736D556D9C3FF0CC96A96CC78078CCB552D9C7FF8664A8A93387FC3996AAB6CE1FF0E6DAAADB387F839B6AAB6C707C1CC92AB498E001E6695569987FF866DAAB4DCF80F8C92AA9331FFF866D4B5B638001CC96AB498E001E669556D9C3FE1CCB555B338001CC92AA499E000E66D556D9C1FC399AD52D98FC7E3369569338080E64B54B663E0F8CCA55ACCE0F8399A55299";
defparam ram_block1a49.mem_init0 = "8FC7E336B52931C001CCDAAADB181E0736D556D8E0007334AAD263C01E324AA96470781CCB555A6703C1CCD2AB49CF80F19B4A94D8F003CCDABA9271FFF1992AA9271FFF8CDA55ACCE02071B6AAB6C700071B6A2A4CE1FE1CC9555B33C00F192D52998F01E3329529B1E00719A555B6703C1C6D2AB49CF81F1925552661FF8736B5693383E0E64ADA9338000E64AAA9338000E64ADA93383E0E64B56B230FF8736D55B661FFC33255524E3FFF19B5256CC7C0F1994A94D8F0078C96AB498F0078C96AB498F0078C96AB498F80F99B5AD6CC7FFE392555A671FF8624A52931C003CC96A96CC3FFC336956931C0038DB5552670FE0E6D2AB6CC3FF8664AAA4CC7F";

cyclonev_ram_block ram_block1a73(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a73_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a73.clk0_core_clock_enable = "ena0";
defparam ram_block1a73.clk0_input_clock_enable = "ena0";
defparam ram_block1a73.clk0_output_clock_enable = "ena0";
defparam ram_block1a73.data_interleave_offset_in_bits = 1;
defparam ram_block1a73.data_interleave_width_in_bits = 1;
defparam ram_block1a73.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a73.init_file_layout = "port_a";
defparam ram_block1a73.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a73.operation_mode = "rom";
defparam ram_block1a73.port_a_address_clear = "none";
defparam ram_block1a73.port_a_address_width = 13;
defparam ram_block1a73.port_a_data_out_clear = "none";
defparam ram_block1a73.port_a_data_out_clock = "clock0";
defparam ram_block1a73.port_a_data_width = 1;
defparam ram_block1a73.port_a_first_address = 24576;
defparam ram_block1a73.port_a_first_bit_number = 1;
defparam ram_block1a73.port_a_last_address = 32767;
defparam ram_block1a73.port_a_logical_ram_depth = 65536;
defparam ram_block1a73.port_a_logical_ram_width = 24;
defparam ram_block1a73.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a73.ram_block_type = "auto";
defparam ram_block1a73.mem_init3 = "03FC03FC03FC01FE00FF803FE007FE003FF8007FFC000FFFFC000003FFFFFFFFFFFFFFFFF800003FFF8007FE00FF00FE07F03E0FC1E0F0787870F1E3871C71C638C6318C663319999999993366CD936C92492496D25A5AD294A56AD52A9555AAAAAAAAAB555AAD52B5294B5A4B49249249B264CD99998CCE739C638F1C3C3C1F03F007FF80000001FFE01FC1F07870E38E39CE673333664D924924B4B4A56AD56AAAAAAAAB55AB5AD2D2DB6D9366CCCCE6318E38F1F0F81FE0003FE0003FC0F87870E718C666664C936D25A5AD5AAD555555AAD4A52DA49364CC9CCC638E3C3C1F801FFFFF801F83C3C71CE63332649B692D6A54AAAAAAA55AD696DB24CCCCCE";
defparam ram_block1a73.mem_init2 = "71C78781FC0000007F03C3C71CC6666CDB6D2D2B55AAAAB55A9696DB26CCC6718F0F07F0000003F83C38E31999936DB4A52A95555AA5296DB66CCC671C783F003FF801F878E39CCCD936D2D4A955552AD696D93666318F1F03FF00FFE0F8F18C666C924B5AB55554A94B49B266739C3C1FC0000FF0F0E3199936DB5AD555554AD2DB664E638E1F00FFFC03E1C71999B2494A554B556A5B6D9999C71E07FFFFF81E1CE7326C9695AAAAAB5ADB6CCCC71C3F000001F871CE664DA4A55AAB55A5B6C99CE387C03FE00F8718CCD925AD52AB54A5B64CC638F03FFFFC0F1C6666496952AAA54B6DB3338E1F000001F0E3999B6DAD52A956B69B3338E1F00000FC38C6";
defparam ram_block1a73.mem_init1 = "64DB4AD5554AD249998E3C1FFFFE0F1C666C96956AB54B4933318F07FFFFC1C3199B2DAD5555296D9339C3C07FF01E18C6CDA5A9554AD6D9339C3C07FE03C39CC9B4B54AB56B6D998E3C0FFF81E18CCDB6956AD52926CC63C1FFFFC1C73336D295554A5B26638F007C01E38CC9B4AD554AD24CCC707E007F0E3193694AAAAD6DB331C3E0003F1C666494AAAAB5B64E63C1FFFE0F19D9B6B5555696CCCE3C0FFC078C66C96A554AD24CCC783FFFC1C7336DAD555696CCCE3C03E01E399924AD552B49998E1F803F0E3336D2AD2AD6C99C707FFF878CCC96B5552964CC71F800FC3999B6B5555A49B18F07FF81C7326D6AAAA5B666387FFFF0E7324B52AD5A4CCC";
defparam ram_block1a73.mem_init0 = "783FFC1E3336DAA52A5B6671E03E03C7336D2A52A5B6631F0000F0C64D2D55529266387FFFE1C66496AAAA5B2630F8003E39992D6AAD6933187E00FC7193695555A499C701FC0718D929555692673C1FFC1E7324B5554A4CCC780003C733694AAD69331C3FFFE1CCC929556B6CCE3C00078E66DAD5529266383FFE1E666D6AAAD24CE3C0003C7324B555692663C0780F199B4AAAB49338F0001E39B252AA96D99C7E01F8E66DA5552D3338FC03F1CCDB52AD49331C1FFC1CE4DAD55293631F001F1CCDA55552498E3FFFE1CCDB52AD69338F0003C7325AD5A964C70FFF8399929554B6CC707FE0E336D6AAD6CCC78000F189B5AAB5B673C0F81E336D2AA96D9C";

cyclonev_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 8191;
defparam ram_block1a1.port_a_logical_ram_depth = 65536;
defparam ram_block1a1.port_a_logical_ram_width = 24;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init3 = "736D2AA96D98F03E079CDB5AAB5B231E0003C666D6AAD6D98E0FFC1C66DA5552933383FFE1C64D2B56B499C78001E3992D6A95B6670FFFF8E32495554B6671F001F18D929556B64E707FF07199256A95B6671F807E399969554B6CCE3F00FC7336D2AA949B38F0001E39925AAAA5B331E03C078CC92D555A499C7800078E6496AAAD6CCCF0FFF838CC929556B6CCE3C00078E66DAD552926670FFFF871992D6AA52D99C780003C6664A5555A499CF07FF079CC92D555293631C07F01C7324B55552D931C7E00FC31992D6AAD693338F8003E18C9B4AAAAD24CC70FFFFC38CC9295556964C61E0001F18CDB4A94A96D99C780F80F1CCDB4A94AB6D998F07FF83C";
defparam ram_block1a1.mem_init2 = "6664B56A95A499CE1FFFFC38CCDB4AAAAD6C99C703FFC1E31B24B5555ADB33387E003F1C664D29555AD26663C3FFFC1C7326D6A96A96D998E1F803F0E33325A9556A493338F00F8078E666D2D5556B6D99C707FFF83C666496A554AD26CC63C07FE078E666D2D5555ADB3731E0FFFF078CE4DB5AAAAA524CCC71F8000F87199B6D6AAAA52D9318E1FC00FC1C666496A5556A5B26638F007C01E38CC9B4A5555296D999C707FFFF078C66C92956AD52DB66630F03FFE078E3336DAD5AA55A5B26738780FFC078739936D6A5552B4B66C630F01FFC078739936D2955556B69B3318707FFFFC1E3199925A55AAD52D26CCC71E0FFFFF078E3332496A55556A5B64C";
defparam ram_block1a1.mem_init1 = "C6387E00001F0E3999B2DAD52A956B6DB3338E1F000001F0E3999B6DA54AAA952D24CCCC71E07FFFF81E38C664DB4A55AA956B49366631C3E00FF807C38E7326DB4B55AAB54A4B64CCE71C3F000001F871C6666DB6B5AAAAAB52D26C99CE70F03FFFFFC0F1C733336DB4AD55A554A5249B3331C70F807FFE01F0E38CE4CDB696A5555556B5B6D933318E1E1FE00007F078739CCC9B25A52A55555AB5A4926CCC631E3E0FFE01FF81F1E318CCD936D2D6A955552A5696D93666738E3C3F003FF801F83C71CC666CDB6D294AB55552A94A5B6D9333318E38783F8000001FC1E1E31CC666C9B6D2D2B55AAAAB55A9696DB66CCCC671C78781FC0000007F03C3C71C";
defparam ram_block1a1.mem_init0 = "E6666649B6D2D6B54AAAAAAA54AD692DB24C9998CE71C78783F003FFFFF003F07878E38C6672664D924B694A56AB5555556AB56B4B496D9264CCCCC631CE1C3C3E07F8000FF8000FF03E1F1E38E318CE6666CD936DB69696B5AB55AAAAAAAAAD56AD4A5A5A49249364CD9999CCE738E38E1C3C1F07F00FFF00000003FFC01F81F0787871E38C739CE6633333664C9B24924925A4B5A5295A956AB555AAAAAAAAAB5552A956AD4A5296B4B496D24924926D9366CD99333333333198CC6318C638C71C71C38F1E1C3C3C1E0F07E0F81FC0FE01FE00FFC003FFF800003FFFFFFFFFFFFFFFFF8000007FFFE0007FFC003FF800FFC00FF803FE00FF007F807F807F80";

cyclonev_ram_block ram_block1a25(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.clk0_output_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "rom";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "clock0";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 8192;
defparam ram_block1a25.port_a_first_bit_number = 1;
defparam ram_block1a25.port_a_last_address = 16383;
defparam ram_block1a25.port_a_logical_ram_depth = 65536;
defparam ram_block1a25.port_a_logical_ram_width = 24;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init3 = "FC664AAA4CC3FF866DAA96CE0FE1CC9555B638007192D52D987FF866D2AD267800719294A48C3FF1CCB554938FFFC66D6B5B33E03E325AAD263C01E325AAD263C01E325AAD263C01E3652A5331E07C66D495B31FFF8E495549987FF0CDB556D9C3FE189AD5A4CE0F83992B6A4CE0003992AAA4CE0003992B6A4CE0F83992D5AD9C3FF0CC9554931F03E725AA96C70781CDB554B31C00F1B2952998F01E332956931E00799B5552670FF0E64A8ADB1C001C6DAAADB1C080E66B54B663FFF1C92AA9331FFF1C92BAB667801E3652A5B31E03E725AA96670781CCB555A6703C1C4D2AA498F0078C96AA599C000E36D556D9C0F031B6AAB667000719295AD98FC7E3";
defparam ram_block1a25.mem_init2 = "32954B3383E0E66B54A663E0F8CDA55A4CE0203992D52D98FC7E336956B3387F0736D556CCE000F324AA9267000399B555A670FF8736D552CCF000E325AAD26700038DB5A56CC3FFF1992AA9263E03E765AAB6CC3FFC332D552CCF000E325AA926707C1C6DAAADB383FC39B6AAB6CE1FF0E6DAAAD3387FC3992A2A4CC3FFC736955A663C03C66D2AD2661FF8736D556D9C3FE1CC95A564E7E1F8CDA552D9C7FFE332D552CCE0003992554B630FFC39B6AAB4CE3FFC732D55699C7FF8E65AAAD330FFF0CC953524E3FFF8CDA556931C001C64B556998F81F19B4AAD333C00F19B4AB5938FFFC736954A6C7000799B5556D8E0F838C94A9499C3FE1CC96AA59987";
defparam ram_block1a25.mem_init1 = "FF0E6DAAA9331F03E332D552CCE1FF0E64A54A4CE1FF0E6695569B9E0078CDA556931C000E324AAA499E000719255524C700038C92AA966703E0E36D6B52661FFF0CC94AD6D8E1FE1C6DAD6A4CC3FFE1992D569330FFF8E65A92B6C60FF87324AAB498E02038D96AAD36380C0F324AAADB387FFC736D555B2307FE1CC94AB5B31E003C66D6AD6D8C1FF0E66D5952663E01E33256B5B670FFF0C4D2AAB6CE3FFF0CC92AAD26383F07192D552D9C7C0F8E6D2AAD26383F07192D556D98F001E3369552D98F000F19252B52661F8FE3325AA96CCE07C0E66D2AB4938F007C66DAAA964E3FFFC736D55526678003C64D6AB5B31C000719B4AA96CCF0380E765AAA92";
defparam ram_block1a25.mem_init0 = "670FFF0E649555A6E703E071925554B231F83F199A5556D99E0003CCCB5552D9C7801E3934AAA5B31E000719B6AAADB31C000F19B6AAADB31C00079D92956B6671FFF87325AAAD2671FFFE3992D5569338FFFF0CC92AAADB31E000F19B6ADAB6CE3C00F8CC96AAB4D9C7FFF8626D6AB5B230FFFF1CC92AAADB33C1FC1C66DAAAA499C7C07C3334AD2A499C3FFF0E6495A95B671E001E3324AAAB6CCE0FFC1CCDB5555B663C00038CDB5AA52CCE3F87E199B5AAB4931C3FFC38C92D55AD9987C07E3992D5552C8C70000E3324AAAB499C7800F0CC92956A4CCE1FFF8633695552C98E1FFF0E664A556B6CC703F03CE4D2A5A964E703FC1E664B55569331E0001E";

cyclonev_ram_block ram_block1a98(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a98_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a98.clk0_core_clock_enable = "ena0";
defparam ram_block1a98.clk0_input_clock_enable = "ena0";
defparam ram_block1a98.clk0_output_clock_enable = "ena0";
defparam ram_block1a98.data_interleave_offset_in_bits = 1;
defparam ram_block1a98.data_interleave_width_in_bits = 1;
defparam ram_block1a98.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a98.init_file_layout = "port_a";
defparam ram_block1a98.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a98.operation_mode = "rom";
defparam ram_block1a98.port_a_address_clear = "none";
defparam ram_block1a98.port_a_address_width = 13;
defparam ram_block1a98.port_a_data_out_clear = "none";
defparam ram_block1a98.port_a_data_out_clock = "clock0";
defparam ram_block1a98.port_a_data_width = 1;
defparam ram_block1a98.port_a_first_address = 32768;
defparam ram_block1a98.port_a_first_bit_number = 2;
defparam ram_block1a98.port_a_last_address = 40959;
defparam ram_block1a98.port_a_logical_ram_depth = 65536;
defparam ram_block1a98.port_a_logical_ram_width = 24;
defparam ram_block1a98.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a98.ram_block_type = "auto";
defparam ram_block1a98.mem_init3 = "070C6326496B56AAB56B69B3331C707F800FF0F1C6666CB6B52AAAD5A5B66CE638781FFFF81F1C73336496B55AA55296D93331C70FC00001F071CE66C925AD555552B492666638E0FE0001FC3C71999B25A52AAAAAD696C9999CE1E0FFFFFF078739899B6D2955AB55296DB26631C783F8001FC1E38CE6CDB694AA556AB5A49326738E1E03FFFF01E1C7333364B4A556AD54A5B6D9999C70F03FFFFF03C38C6666DB694AA554AB5A5B66CCE71C3E03FFFE03E1C7319B36D252AD555AA52DB64CCE73C7C1FFFFFF03C38C6666C92D2B555555294924D998C71E1FC00000FC1E38CE66C924A52AB54AAD4B69B266631C3C1FE0003FC1E1CE3333649694A95555AB";
defparam ram_block1a98.mem_init2 = "5A5B64CCCE71C3E07FFFFF01E1E318CCD92496B54AAAAD5AD6DB66CCE738787E0000003F0F1C733B326DA5AD5AAAAAD5AD2493666739E3C3F8000001F878718CCCC9B6D2D6AB5556AB5A5B6D9B319CE1C3E01FFFFF01F0F1C6333326DB4B52AD5556AB5A5B6D9B3398E38F83F800001FC1F1C718CCC9924B4B52AA96AAB5296D26CD99CC71C783F80000007E0F0E39CCCCC9B6DA52954AAAA55294B6DB664CE639C3C3E01FFFFFE03E0E1C731999B26D25A56A955556AB5AD25926CCCCE71C70F81FF00003FE07C38E39CCCCC9B6DA5A56AB55556AB5296D26D9B3319CE38787E01FFFFFF80FC3C38E739999B26DB4B5AD52AAAAAB54AD2D249366CCE631C71E";
defparam ram_block1a98.mem_init1 = "1F81FFE003FFC07C3C38E739999936496D2D6AD54AAAA556AD696D24D93333318C71E1E0FC03FFFFFF007E0F0E38E3399999364925A5295AA955556AA54A52DA49B66CCCCC631C71E1F07F000FFFE001FC1F0F1E31CE6333264D924B694A56AB55555552A95AD2D25B64D93333398C71C78783E03FF000000FFC07E1F1E3C639CC66664C9B2496D2D6B52AD555555554AB5294B496DB24C9993999CE71C70E1E0FC0FF8000000007FC0FC3E1E38E38C6733333366C924925A5AD6A55AAA555555AAA54AD4A5A5B6936D9326666667318E31E38787C1F01FF0000FFF80007F80FC1F0F1E38738C6339999999326C936D24B4B4A52B54AA55552AA95554AA54A94";
defparam ram_block1a98.mem_init0 = "A5A5A5B6DB6D9366CC99998CC6739C71C71E3C3E1F03F01FE000FFFFFFFFC003FE01F83E0F070F1E38E39C63398CCCE6CCCD993649B6DB6DA4B4B4A5AD4AD5AA556AAA95555554AAAB552AD52B5A94B5A5A4B4924B64936C9B366CCD999998CCE6739CE718E38E3871E1C3C3E1F07C0FC07F007FE000FFFFFFFFFFFFFFFE000FFC01FE03F03F07C1F0F87878F0E1C78E38E38E71CE739CE73198CCE6666333266666CCD9B366C9936C9B64936DB6DB6DB492DB49692D2D2D2D29694A5AD6B5295A95A95AB56AD5AA552AD54AAD55AAAD554AAAB55555AAAAAAA9555555555555555555555554AAAAAAAA9555555AAAAAB55554AAAA95554AAAA55552AAAD5552";

cyclonev_ram_block ram_block1a122(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a122_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a122.clk0_core_clock_enable = "ena0";
defparam ram_block1a122.clk0_input_clock_enable = "ena0";
defparam ram_block1a122.clk0_output_clock_enable = "ena0";
defparam ram_block1a122.data_interleave_offset_in_bits = 1;
defparam ram_block1a122.data_interleave_width_in_bits = 1;
defparam ram_block1a122.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a122.init_file_layout = "port_a";
defparam ram_block1a122.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a122.operation_mode = "rom";
defparam ram_block1a122.port_a_address_clear = "none";
defparam ram_block1a122.port_a_address_width = 13;
defparam ram_block1a122.port_a_data_out_clear = "none";
defparam ram_block1a122.port_a_data_out_clock = "clock0";
defparam ram_block1a122.port_a_data_width = 1;
defparam ram_block1a122.port_a_first_address = 40960;
defparam ram_block1a122.port_a_first_bit_number = 2;
defparam ram_block1a122.port_a_last_address = 49151;
defparam ram_block1a122.port_a_logical_ram_depth = 65536;
defparam ram_block1a122.port_a_logical_ram_width = 24;
defparam ram_block1a122.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a122.ram_block_type = "auto";
defparam ram_block1a122.mem_init3 = "00F0E7364B5AAAB5A4CCC71F8003E1C664DAD5A956926673C1FFFE0F399925AB56A96D998E3F0003E1CE6C9295554A593318780000F8E666DA555552DB3338F0000078E666DAD5555ADB3338780000F0C6649295554A49339C3E0003E1CC4C96A5552B6D998E1F800FC38CCDB4AD55A96C99CE1FC01FC38CCDB4AD55A96D998E3F0003E1CE649295555ADB2738E03FF81E319B6D2AAAAD6D999C3C00007873336D6AAAA96DB318F07FFE0F1CCD92D5AAD4B4D98C780FFC0F1CCCDA5AAAA94936738780003E38CC9A5AAAAA524CCC787FFFF07199925A9552B49B318F03FF81E39C9B6B55556B6CCCE3C0FFC078C66C96A555A96C99C70FE03FC38CCD96955552";
defparam ram_block1a122.mem_init2 = "D2666387E003F0E33325A55554B49998E1F800FC38CCD96B55552D2666387C001F8739924B56A952DB3338F01FE03C319B25AD554AD26CC71E03F8078E666DA54AA54B64CC71F00003E39CD9252AAAA524D8CE1F0000F8739924B54AD52DB3338F03FF80E18CD92D4AAA56936631E07FFC0F18CD92D4AAAD6926671E0FFFF071CCCDA5AAAAA5A4CCC70F8001F873993695AAAD4B6CCC71F00003E18CCDB6B5555AD26CC71E07FE03C73136DA9555A96C99CE1F0000F873993694AAAB5A4D98C783FFFC1E399924A55556B49919C7807F00F1CE4C9695555296CCCC787FFFFC3CE6649295555ADB66671F01FC03C719934B52AA54B6CCCE3C0FFF81E3999B694A";
defparam ram_block1a122.mem_init1 = "AAB5A4D98C787FFFF878C64DB4A5556A5B66671E07FFE0F1C66C92955554B49999C7C07FC078E736496AD54A96D9318E1FC00FE1C6326DA56AA95A593338F07FFFC1E39993695AAAD5B4D998E1F00007C38CCC92D6AAAB5A4D99CF1F8001F8718C9B6952AA56B6CCCC707E003F8718CDB6D4AAAA52D93318783FFF81E3999B6D2AB6AB5B6CCC63C0FFFE0F0C666DA5AAAAAD2DB3318F03FFFC1E38CC924AD5556B4936338F01FFE03C739B2494AAAAB5B6C98C70FE001FC38C66C96955555ADB66671C3FE07F838E666DA52AAAA52DB3339E1F8003F0F3999B6D6AAAAB5A4D99C71F00000F8F399B25A55AB54A493331C7807FE03C7199934B56AAD5A5B26738";
defparam ram_block1a122.mem_init0 = "F03FFFC0F1CE64DA5A9554AD6D9331C707FFFF83C73993696AD55AB4B64CC71C1FFFFF838E736492952A95696C998C787F803FC3C63326D2D52AB56B6D999C70F80001F8719CD925AD5555296D9339C783FFFFC1E38CCD96D6AB5AAD69366638E0FFFFFC1E39CD9B695AAAAB5A5933318783FFFFC1E39CCD92D2A5552A5A4D99CE3C1FFFFF078E3336496A55556A5B6CCCE78F800C0078718CC9B4B52AAAD4B49B331C707F001FE1E3199924B5AAAAAD6924CCCE387E0000FE1C73332496B55555296D93338E3E01FF8078718CC9B694AAAAA94B6D999CE1E07FFFE078E319B2496A55556A5A49999CE1F01FFF01F1C73336DB5AB5552A5A49B339C783FC00FF";

cyclonev_ram_block ram_block1a146(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a146_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a146.clk0_core_clock_enable = "ena0";
defparam ram_block1a146.clk0_input_clock_enable = "ena0";
defparam ram_block1a146.clk0_output_clock_enable = "ena0";
defparam ram_block1a146.data_interleave_offset_in_bits = 1;
defparam ram_block1a146.data_interleave_width_in_bits = 1;
defparam ram_block1a146.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a146.init_file_layout = "port_a";
defparam ram_block1a146.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a146.operation_mode = "rom";
defparam ram_block1a146.port_a_address_clear = "none";
defparam ram_block1a146.port_a_address_width = 13;
defparam ram_block1a146.port_a_data_out_clear = "none";
defparam ram_block1a146.port_a_data_out_clock = "clock0";
defparam ram_block1a146.port_a_data_width = 1;
defparam ram_block1a146.port_a_first_address = 49152;
defparam ram_block1a146.port_a_first_bit_number = 2;
defparam ram_block1a146.port_a_last_address = 57343;
defparam ram_block1a146.port_a_logical_ram_depth = 65536;
defparam ram_block1a146.port_a_logical_ram_width = 24;
defparam ram_block1a146.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a146.ram_block_type = "auto";
defparam ram_block1a146.mem_init3 = "FE007F83C7399B24B4A9555AB5B6D999C71F01FFF01F0E733324B4AD5554AD249B318E3C0FFFFC0F0E73336DA52AAAAA52DB26631C3C03FF00F8E399936D2955555AD249999C70FE0000FC38E666492D6AAAAB5A4933318F0FF001FC1C7199B25A56AAA95A5B26631C3C006003E3CE666DB4AD5554AD24D998E3C1FFFFF078E73364B4A9554A969366738F07FFFF83C3199934B5AAAAB52DB36738F07FFFFE0E38CCD92D6AB5AAD6D366638F07FFFF83C739936D2955556B4936731C3F00003E1C73336DAD5AA95696C998C787F803FC3C63326D2D52A952924D9CE383FFFFF071C664DA5AB556AD2D9339C783FFFFC1C719936D6A5552B4B64CE71E07FFF81E";
defparam ram_block1a146.mem_init2 = "39CC9B4B56AAD5A593331C780FFC03C7199924A55AB54B49B339E3E00001F1C73364B5AAAAAD6DB3339E1F8003F0F3999B694AAAA94B6CCCE383FC0FF871CCCDB6B555552D26CC6387F000FE1C6326DB5AAAAA5249B39C780FFF01E398D925AD5556A4926638F07FFF81E3199B696AAAAB4B6CCC61E0FFFE078C666DB5AADAA96DB3338F03FFF83C31993694AAAA56DB6631C3F800FC1C6666DAD4AA952DB2631C3F0003F1E73364B5AAAAD692666387C0001F0E33365B56AAB52D93338F07FFFC1E399934B52AAD4B6C98C70FE007F0E31936D2A556AD24D9CE3C07FC07C733325A555552926CC71E0FFFC0F1CCCDB4AD554A5B64C63C3FFFFC3C63364B5AAA";
defparam ram_block1a146.mem_init1 = "A52DB3338F03FFE078E666DA54AA95A59331C7807F01F1CCCDB6B55552924CCE787FFFFC3C6666D2955552D264E71E01FC03C731325AD5554A493338F07FFF83C63364B5AAAA52D9339C3E0001F0E7326D2B5552B6D919C780FFC0F1C66C96B5555ADB66630F80001F1C666DA56AAB52D9339C3F0003E1C6664B4AAAAB4B66671C1FFFE0F1CCC92D6AAA56936631E07FFC0F18CD92D4AAA56936630E03FF81E3999B6956A55A49339C3E0001F0E636494AAAA94936738F80001F1C664DA54AA54B6CCCE3C03F80F1C66C96A5556B49B318780FF01E3999B6952AD5A49339C3F0007C38CCC9695555AD3666387E003F0E33325A55554B49998E1F800FC38CCC96";
defparam ram_block1a146.mem_init0 = "955552D3666387F80FE1C7326D2B554AD26CC63C07FE078E666DAD5555ADB2738F03FF81E319B25A9552B493331C1FFFFC3C666494AAAAB4B26638F80003C39CD9252AAAB4B66671E07FE03C63365A56AB56936671E0FFFC1E319B6D2AAAAD6D999C3C00007873336D6AAAA96DB318F03FF80E39C9B6B55552924CE70F8001F8E3336D2B556A5B666387F007F0E7326D2B556A5B666387E003F0E3336DA9554AD264670F8000F8739924A55552924CC61E00003C3999B6B55556B6CCCE3C00001E3999B6955554B6CCCE3E00003C319934A55552926CE70F8001F8E3336D2AD5AB493339E0FFFF079CCC92D52B56B64CC70F8003F1C6664B5AAAB5A4D9CE1E00";

cyclonev_ram_block ram_block1a170(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a170_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a170.clk0_core_clock_enable = "ena0";
defparam ram_block1a170.clk0_input_clock_enable = "ena0";
defparam ram_block1a170.clk0_output_clock_enable = "ena0";
defparam ram_block1a170.data_interleave_offset_in_bits = 1;
defparam ram_block1a170.data_interleave_width_in_bits = 1;
defparam ram_block1a170.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a170.init_file_layout = "port_a";
defparam ram_block1a170.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a170.operation_mode = "rom";
defparam ram_block1a170.port_a_address_clear = "none";
defparam ram_block1a170.port_a_address_width = 13;
defparam ram_block1a170.port_a_data_out_clear = "none";
defparam ram_block1a170.port_a_data_out_clock = "clock0";
defparam ram_block1a170.port_a_data_width = 1;
defparam ram_block1a170.port_a_first_address = 57344;
defparam ram_block1a170.port_a_first_bit_number = 2;
defparam ram_block1a170.port_a_last_address = 65535;
defparam ram_block1a170.port_a_logical_ram_depth = 65536;
defparam ram_block1a170.port_a_logical_ram_width = 24;
defparam ram_block1a170.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a170.ram_block_type = "auto";
defparam ram_block1a170.mem_init3 = "95556AAA95554AAAA55552AAAA55555AAAAAB5555552AAAAAAAA5555555555555555555555552AAAAAAB55555AAAA5556AAB556AA556A954AB56AD5AB52B52B5295AD6B4A52D29696969692D25B6925B6DB6DB6D924DB26D9326CD9B3666CCCCC9998CCCCE663319CE739CE71CE38E38E3C70E1E3C3C3E1F07C1F81F80FF007FE000FFFFFFFFFFFFFFFE000FFC01FC07E07C1F0F87870F1C38E38E31CE739CCE66333333666CD9B26D924DA4925A4B4B5A52B5A956A955AAAA55555552AAAD54AB56A56B4A5A5A4B6DB6DB24D9336666CE6663398C738E38F1E1C1E0F83F00FF8007FFFFFFFE000FF01F81F0F878F1C71C739CC663333266CD936DB6DB4B4B4A";
defparam ram_block1a170.mem_init2 = "52A54AA55552AA95554AA55A94A5A5A496D926C99333333398C639C38F1E1F07E03FC0003FFE0001FF01F07C3C38F18E319CCCCCCC9936D92DB4B4A56A54AAB555554AAB54AD6B4B4924926CD999999CC638E38F0F87E07FC000000003FE07E0F0E1C71CE73339332649B6D25A5295AA5555555556A95AD696D249B264CCCC6738C78F1F0FC07FE000001FF80F83C3C71C63399999364DB49696B52A95555555AAD4A52DA49364C9998CE718F1E1F07F000FFFE001FC1F0F1C718C66666CDB24B694A54AAD55552AB5294B4924D93333398E38E1E0FC01FFFFFF807E0F0F1C6319999936496D2D6AD54AAAA556AD696D24D9333339CE38787C07FF800FFF03F0";
defparam ram_block1a170.mem_init1 = "F1C718CE66CD9249696A55AAAAAA956B5A5B6C9B33339CE38787E03FFFFFF00FC3C38E73199B36C96D295AAD5555AAD4B4B6DB26666738E387C0FF80001FF03E1C71CE6666C93496B5AAD55552AD4B496C9B33319C70E0F80FFFFFF00F878738CE64CDB6DA52954AAAA55294B6DB26666738E1E0FC0000003F83C71C673366C96D295AAAD2AA95A5A493266631C71F07F000003F83E38E3399B36DB4B5AAD5556A95A5B6C99998C71E1F01FFFFF00F870E7319B36DB4B5AAD555AAD696DB2666631C3C3F0000003F878F39CCCD92496B56AAAAB56B4B6C99B99C71E1F8000000FC3C39CE66CDB6D6B56AAAA55AD2493666318F0F01FFFFFC0F871CE6664DB4B5";
defparam ram_block1a170.mem_init0 = "AB55552A52D24D9998E70F07F8000FF078718CCC9B2DA56AA55AA94A4926CCE638F07E000007F0F1C63336492529555555A96926CCCC638781FFFFFF07C79CE664DB694AB5556A9496D9B319C70F80FFFF80F871CE66CDB4B5AA554AA52DB6CCCC638781FFFFF81E1C733336DB4A556AD54A5A4D9999C70F01FFFF80F0E39CC9924B5AAD54AA52DB66CE638F07F0003F83C718CC9B6D2955AB55296DB32339C3C1FFFFFE0F0E733326D2D6AAAAA94B49B3331C787F0000FE0E38CCCC925A9555556B4926CCE71C1F000007E1C7199936D2954AB55AD24D999C71F03FFFF03C38CE6CDB4B56AAA95ADA6CCCC71E1FE003FC1C71999B2DAD5AAAD5AD24C98C61C1";

cyclonev_ram_block ram_block1a50(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a50_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a50.clk0_core_clock_enable = "ena0";
defparam ram_block1a50.clk0_input_clock_enable = "ena0";
defparam ram_block1a50.clk0_output_clock_enable = "ena0";
defparam ram_block1a50.data_interleave_offset_in_bits = 1;
defparam ram_block1a50.data_interleave_width_in_bits = 1;
defparam ram_block1a50.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a50.init_file_layout = "port_a";
defparam ram_block1a50.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a50.operation_mode = "rom";
defparam ram_block1a50.port_a_address_clear = "none";
defparam ram_block1a50.port_a_address_width = 13;
defparam ram_block1a50.port_a_data_out_clear = "none";
defparam ram_block1a50.port_a_data_out_clock = "clock0";
defparam ram_block1a50.port_a_data_width = 1;
defparam ram_block1a50.port_a_first_address = 16384;
defparam ram_block1a50.port_a_first_bit_number = 2;
defparam ram_block1a50.port_a_last_address = 24575;
defparam ram_block1a50.port_a_logical_ram_depth = 65536;
defparam ram_block1a50.port_a_logical_ram_width = 24;
defparam ram_block1a50.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a50.ram_block_type = "auto";
defparam ram_block1a50.mem_init3 = "0FFFF01E1CE666C9695AAAAB5ADB66C671C1F80001F871CE66C9694AAAAA56924CCCE387C00000F878CE64DB4B54AA95296C9999C787E0001F838E6664DA52A952A96926CCE71E07FFFF81E39CCD925A556955AD24D98C71E07FFF80F1C6666DB4A55555AD249999C787F000FE0E39CD9B694AAAAAD69264E6387803F807C38CCCDB695AAAAD4B6D9998E1F000001F1C6336492955555292C999CE1E01FF80F8E33B36DA54AAA54B6D9998E1E000003E1CE664DA52AAAAB5A4D998C783FFFFE0F1CE64DA5A95552B49266638F01FFF81E38CCC925A9555AB49266638F80FFC07C7199934B52AAA56924CCC70F007C01F1C6666DA56AAAB5A593331C3E00001F0";
defparam ram_block1a50.mem_init2 = "E3332696B5554AD24999C70FC0007E1C6336496AD556A5A4CCCE383FFFFF071CCCDB6956AB56B6C998E3C1FFFF078E3326D2D54955A5B36738F01FFE03C7199B6D2A554A96DB3318F03FFFC0F18CCDB6B54AD52924CCE70FC0003F0E73324B4AAAAA5249998E3E00001F1C6366D2D5AA55A5B3731C3E00007C718C9B6952AA54B6C99CE1F00001F1C666492955556B6D999C781FFFC0E18CC9A4AD555A96C999C783FFFF071CE4D96B55554B49B318F0FFFFF878CE4DB6A5555A924D9CE1E00000F0E636492B5554A5B66671E07FFE078E666DA56AAA5692666387E0007E1CE66DB4A955A969B331C3E0000F873993694AAAA52DB33187807E01E1CCCDB6B555";
defparam ram_block1a50.mem_init1 = "5696D99CE1F00007C39CC9B4AD555A924CCC70FC001F8F399B6D6AAAA94936638F01FF81E18CC925AA56A969B339C3F0007E1CE66DB4AAAAA524C8CE1E00001E18CCD96B55552964CCE783FFFF079CCC9252AAAB5B6CCC70F8000F87199B2D2AAAAD6DB338E1FF0FF0718D9B4A55552924CCE383FFFF0F18CDB6952AD5A59331C7C000078731325AD5556B4D998E3E0000F8E3336DAD5556B6D998E3F0001F0E3326D2B554AD24CCE787FFFF871CCD96952A55A49998F0FFFFF8718D924AD554A5B267387E001F87199B6D6AAAB5A6CCC70F8001F0E3336D2B555AD24CCE383FFFC1E319B6D2A92A96DB318F07FFF078C66DB4AB5AA5A6CC63C1FFFC1E399B2D";
defparam ram_block1a50.mem_init0 = "2A92A96D9318F03FFE0F1CCC9252AAAD6DB331C7E0007C38CC9B4A954A96D998E3F0001F0C666CB5AAAB5A4998C7C07F01E38CD96D5AA95A49998E0FFFFE1E33324A55555A49339C3E0007E38CCDB6A5552B6D919C3E0001F0E666DA56AA54B64CE787F01FC3CE64D254AAD4B6CCC71F0001F8E3326D6AD4AB493331E1FFFF838C64DA52AAA52D9B98F07FFF078CCCDA52AAA52D9B98F07FFF078C64DB5AAAAD6DB338E1FFFFC3C666494AAAAB493631C3FC0FE1E732692A552A5B267387F007F0E7326D2A552A5B267387F80FE1C636496AAAA9493339E0FFFF838C64DA56AA95A4D98E3C00003C719B25A9556A493331E0FFFF071CCDB6955552D26663C3FF";

cyclonev_ram_block ram_block1a74(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a74_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a74.clk0_core_clock_enable = "ena0";
defparam ram_block1a74.clk0_input_clock_enable = "ena0";
defparam ram_block1a74.clk0_output_clock_enable = "ena0";
defparam ram_block1a74.data_interleave_offset_in_bits = 1;
defparam ram_block1a74.data_interleave_width_in_bits = 1;
defparam ram_block1a74.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a74.init_file_layout = "port_a";
defparam ram_block1a74.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a74.operation_mode = "rom";
defparam ram_block1a74.port_a_address_clear = "none";
defparam ram_block1a74.port_a_address_width = 13;
defparam ram_block1a74.port_a_data_out_clear = "none";
defparam ram_block1a74.port_a_data_out_clock = "clock0";
defparam ram_block1a74.port_a_data_width = 1;
defparam ram_block1a74.port_a_first_address = 24576;
defparam ram_block1a74.port_a_first_bit_number = 2;
defparam ram_block1a74.port_a_last_address = 32767;
defparam ram_block1a74.port_a_logical_ram_depth = 65536;
defparam ram_block1a74.port_a_logical_ram_width = 24;
defparam ram_block1a74.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a74.ram_block_type = "auto";
defparam ram_block1a74.mem_init3 = "AAA95556AAA95554AAAAD5554AAAAB555552AAAAA955555556AAAAAAAAAAAAAAAAAAAAAAAAAAAA95555552AAAA5555AAAD556AA554AA552AD52A54A952B52B5295AD6B5AD296B4B4B4B4B496D25B4925B6DB6DB24936C9B64D93264C99B333666666666733399CCE7318C739C738E38E3871E3C3878783C1F07C1F80FC03FC00FFF000007FFFFFFE00001FFE007F80FC0FC1F0783C3C7871E38E38C738C673198CCCCCCCCD99326C9B64924925B49696B4A52B52A55AAD554AAAAAAAAA9555AAD52A52B5AD2D2D25B6DB6C9364C99B33333399CC631C638F1C3C7C3C1F81FC03FF80000000001FFC03F81F07C3C3871C71CE7398CCCCCCC99364DB6DB6969694";
defparam ram_block1a74.mem_init2 = "A56AD52AA95555552AA956AD4A52D2DA49249B66CC99998CC6718E38E1C3C1F07F00FFF0000003FFC03F03E1E1E38E38C633199993364DB6DB49694A56AD55AAAAAAAB552A56B5A5B49249B264CCCCE6318E38F1E1F07F00FFFF00FFFF00FE0F878F1C739CC66666CD926D24B4A52956AA95555AAA55A94B4B6DB6C9B3333339CE38E1C1E07E00FFFFFFFC01F81E1E3C718C6672664C92492D2D6A54AAAAAAAAB54A5296DA4DB366666739C71C3C3F03FF000001FF81F07871C7399CCD9936DB6D294AD56AAAAAA552B5A5B49364C998CC638E3C3E07F00000000FE07878718E6333366DB6DA5AD4AA555554AA56B4B6DB64C998CE71870F07E00FFFFF003F07";
defparam ram_block1a74.mem_init1 = "871C731999936492D2D4A95555555AB52D25B24CD98CC738F0F07F00000001FC1E1C31CE66664DB6DA52956AAAAAB54A525B6C9B3339CE38F07C03FFFFFC03E0F1C7398CD9B2492D2B56AAAAAB54A5A4924CD9CCE71E3C1FC0000001F83C38E31999936DB4B52A555554A95A5B6D9B3339CE3C3C0FFE007FF03E1C718CCCC9B6DA5A954AAA954AD2D24D99998C71C1E03FFFFFF01E1E38C66664DB696B56AAAAAD5AD25B26CCC631C3C3F8000001F83C71CE6664DB696B56AAAAB56B4B6D9B3318C78781FF803FF03C38E331B36492D6A5555552A5A5B26CCCE71C3C0FF800FFC1E1C73999936D252A555554AD6924D9999C71E1F8000000F83C739CC9936969";
defparam ram_block1a74.mem_init0 = "52AAAAB5696DB66CE638E1F01FFFFC07C38E339B36DB4A55AAAA55AD249B33318E1E07FFFFFE078718CCCC924B5AAD556A94B49B266318F0F801FF007E1C71999936D295AAAAAD4A4B64CCCE71E0FC00001F83C7399993696952AAA95296DB266318F0FC000001F0F1CE664DB694A95552A52DB64CCE71E1F800001F878E73336496B56AAA95296D933318E1E03FFFF01E1C733326DA52A5554A9496C9998E387C01FE00F871C66649A5AD56A954A5B6C99CC70F03FFFFE0F8E3199B25B5AA554AB5A4933331C781FFFFFE0F1C63364DA52A5556AD69364C671C3F000003E1E319992496A55555A96DB26631C3C07FFF01F1C63326DB5A95554A96DB66671C7C";

cyclonev_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 8191;
defparam ram_block1a2.port_a_logical_ram_depth = 65536;
defparam ram_block1a2.port_a_logical_ram_width = 24;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init3 = "7C71CCCDB6D2A55552B5B6C998C71F01FFFC078718CC9B6D2B55554AD24933318F0F800001F871CC64D92D6AD554A94B64D98C71E0FFFFFF03C71999924B5AA554AB5B49B3318E3E0FFFFF81E1C67326DB4A552AD56B4B24CCC71C3E00FF007C38E33326D252A5554A94B6C9999C70F01FFFF80F0E3199936D2952AAAD5AD24D999CE3C3F000003F0F1CE664DB694A95552A52DB64CCE71E1F0000007E1E318CC9B6D2952AAA952D2D933339C783F000007E0F1CE6664DA4A56AAAAB5296D933331C70FC01FF003E1E318CC9B25A52AD556AB5A492666631C3C0FFFFFFC0F0E31999B2496B54AAAB54A5B6D9B398E387C07FFFF01F0E38CE6CDB6D2D5AAAAA95";
defparam ram_block1a2.mem_init2 = "2D2D9326739C783E0000003F0F1C733336492D6A555554A9496D933339C70F07FE003FE07871CE666C9B4B4A9555554AD6924D9B198E38781FF803FF03C3C63199B36DA5AD5AAAAAD5AD2DB64CCCE71C783F0000003F878718C666C9B496B56AAAAAD5AD2DB64CCCC638F0F01FFFFFF80F071C633333649696A552AAA552B4B6DB2666631C70F81FFC00FFE07878E73999B36DB4B52A555554A95A5B6D9333318E38783F00000007F078F1CE673664924B4A55AAAAAAD5A969249B366339C71E0F807FFFFF807C1E38E73999B26DB494A55AAAAAAD5294B6DB64CCCCE71870F07F00000001FC1E1E39C66336649B49695AB55555552A5696924D9333319C71C3";
defparam ram_block1a2.mem_init1 = "C1F801FFFFE00FC1E1C31CE633264DB6DA5AD4AA555554AA56B4B6DB6CD9998CE31C3C3C0FE00000001FC0F878E38C6633264D925B4B5A954AAAAAAD56A5296DB6D933667339C71C3C1F03FF000001FF81F87871C739CCCCCD9B64B6D294A55AAAAAAAAA54AD6969249264CC9CCC631C78F0F03F007FFFFFFE00FC0F070E38E73999999B26DB6DA5A52B54AAB55552AAD5294A5A496C9366CCCCC6739C71E3C3E0FE01FFFE01FFFE01FC1F0F1E38E318CE66664C9B24925B4B5AD4A955AAAAAAAB556AD4A52D25B6DB64D993333198C638E38F0F0F81F807FF8000001FFE01FC1F07870E38E31CC663333266CDB24924B69694A56AD52AA95555552AA956AD4A";
defparam ram_block1a2.mem_init0 = "52D2D2DB6DB64D9326666666339CE71C71C38787C1F03F807FF00000000003FF807F03F0787C7871E38C718C6733999999B3264D926DB6DB4969696B5A94A956AB5552AAAAAAAAA5556AB54A95A94A5AD2D25B4924924DB26C99336666666663319CC639C638E38F1C3C78783C1F07E07E03FC00FFF00000FFFFFFFC00001FFE007F807E03F07C1F0783C3C3878F1C38E38E39C739C6319CE6733999CCCCCCCCCD999B3264C99364DB26D9249B6DB6DB4925B496D25A5A5A5A5AD296B5AD6B5295A95A952A54A956A954AA554AAD556AAB5554AAAA95555552AAAAAAAAAAAAAAAAAAAAAAAAAAAAD55555552AAAAA955555AAAAA55556AAAA55552AAAD5552AAA";

cyclonev_ram_block ram_block1a26(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.clk0_output_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "rom";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "clock0";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 8192;
defparam ram_block1a26.port_a_first_bit_number = 2;
defparam ram_block1a26.port_a_last_address = 16383;
defparam ram_block1a26.port_a_logical_ram_depth = 65536;
defparam ram_block1a26.port_a_logical_ram_width = 24;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init3 = "FF878CCC96955552DB6671C1FFFE0F199924AD552B49B31C78000078E3364B52AAD4B64C6383FFFE0F3999252AAAAD24D8C70FE03FC39CC9B4A954A96C99CE1FC01FC39CC9B4A954A92C99CF0FE07F8718D925AAAAA524CCC787FFFF0E399B6D6AAAB5B64C63C1FFFC1E33B3694AAA94B66663C1FFFC1E33B3694AAA94B64C6383FFFF0F199925AA56AD6C998E3F0001F1C666DA56AA54964CE787F01FC3CE64DA54AAD4B6CCCE1F0000F873136DA9554ADB66638FC000F8739924B55554A49998F0FFFFE0E33324B52AB56D36638F01FC07C63324B5AAAB5A6CCC61F0001F8E3336D2A552A5B266387C000FC7199B6D6AAA94926671E0FFF81E31936D2A92A9";
defparam ram_block1a26.mem_init2 = "69B338F07FFF078C66CB4AB5AA5B6CC63C1FFFC1E319B6D2A92A96DB318F07FFF838E66496B555A96D998E1F0003E1C666CB5AAAAD6DB331C3F000FC39CC9B4A5556A493631C3FFFFE1E33324B54A952D36671C3FFFFC3CE66496A555A96C998E1F0001F8E3336DAD5556B6D998E3E0000F8E33365AD5556B49919C3C00007C719934B56A952DB6631E1FFFF838E6649295554A5B3631C1FE1FF0E399B6D6AAAA969B331C3E0003E1C666DB5AAAA94926673C1FFFF83CE664D295555AD366630F00000F0E626494AAAAA5B6CCE70FC001F87399B2D2AD4AB4926630F03FF01E38CD9252AAAAD6DB339E3F0007E1C666492B5556A5B267387C0001F0E7336D2D5";
defparam ram_block1a26.mem_init1 = "555ADB66670F00FC03C3199B694AAAA52D9339C3E0000F87199B2D2B552A5B6CCE70FC000FC38CCC92D4AAAD4B6CCCE3C0FFFC0F1CCCDB4A5555A924D8CE1E00000F0E736492B5554ADB64E63C3FFFFE1E319B25A55555AD364E71C1FFFF83C73326D2B5556A4B26630E07FFF03C73336DAD55552924CCC71F00001F0E7326DA54AA952DB2631C7C0000F8719D9B4B54AB5696CD8C71F00000F8E3332494AAAAA5A4999CE1F80007E1CE66492956A55ADB66631E07FFF81E3199B6D2A554A96DB331C780FFF01E39CD9B4B55255696C998E3C1FFFF078E3326DAD5AAD52DB66671C1FFFFF838E6664B4AD556AD24D98C70FC0007E1C7332496A5555AD2C9998E";
defparam ram_block1a26.mem_init0 = "1F00000F87199934B5AAAAD4B6CCCC71F007C01E1C666492D4AAA95A593331C7C07FE03E38CCC925AB5552B49266638F03FFF01E38CCC925A95552B4B64CE71E0FFFFF83C633364B5AAAAA94B64CCE70F800000F0E33336DA54AAA54B6D9B98E3E03FF00F0E73326929555552924D98C71F000001F0E33336DA56AAAB52DB6666387C03F803C38CE4C92D6AAAAA52DB36738E0FE001FC3C73332496B55554A5B6CCCC71E03FFFC0F1C6336496B552D54B49366738F03FFFFC0F1CE66C92D2A952A94B64CCCE383F0000FC3C733326D2952AA55A5B64CE63C3E000007C38E666492D4AAAAA52D26CCE71C3F00003F071CC6CDB6B5AAAAB52D26CCCE70F01FFFE0";

cyclonev_ram_block ram_block1a99(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a99_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a99.clk0_core_clock_enable = "ena0";
defparam ram_block1a99.clk0_input_clock_enable = "ena0";
defparam ram_block1a99.clk0_output_clock_enable = "ena0";
defparam ram_block1a99.data_interleave_offset_in_bits = 1;
defparam ram_block1a99.data_interleave_width_in_bits = 1;
defparam ram_block1a99.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a99.init_file_layout = "port_a";
defparam ram_block1a99.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a99.operation_mode = "rom";
defparam ram_block1a99.port_a_address_clear = "none";
defparam ram_block1a99.port_a_address_width = 13;
defparam ram_block1a99.port_a_data_out_clear = "none";
defparam ram_block1a99.port_a_data_out_clock = "clock0";
defparam ram_block1a99.port_a_data_width = 1;
defparam ram_block1a99.port_a_first_address = 32768;
defparam ram_block1a99.port_a_first_bit_number = 3;
defparam ram_block1a99.port_a_last_address = 40959;
defparam ram_block1a99.port_a_logical_ram_depth = 65536;
defparam ram_block1a99.port_a_logical_ram_width = 24;
defparam ram_block1a99.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a99.ram_block_type = "auto";
defparam ram_block1a99.mem_init3 = "55A94A4B6DB264CCC6738E3C3C1F807FFFFFF00FC1E1E38E731999B36C92DA52952AB55552AA56A5A5B6DB266CC66318E1C3C1F80FFFFFFFF00FC1E1C71C633333366DB6D2D295AA55555556A95AD2D249364CCCCCE718F1E1E0FE00FFFFFF007F0787871CE733993364DB692D6B52A95555556AB5294B6924D933667339C71C387C0FE003FFFF001FC0F0F0E38C63319B326C924B4B4AD5AA955555AA95294B4B6DB26CC998CC639C78F0F81FC003FFFE001FC0F078F1CE319CCCC9936492DA5AD6AD54AAAAAA556AD6B4B49249B2666666318E38E1E0F81FE000000003FE07C1E1C71C63198CD99B26DB692D294A954AAAAAAA954A94A5A5B6DB26CD9999CC";
defparam ram_block1a99.mem_init2 = "639C78F0F07E03FF800000FFE01F07C3C71C718CC66664C9B2492DA5AD6AD52AAAAAAAAA55A95A525B4936C993333319CE38E38787C1FC03FFFFFFFFF807F07C3C3871CE3198CCCD9936C924B694B5AB56AAB55555AAA55A94A5A5B4926D9B366667339C638E1C3C1F03F003FFFFFFFFC00FC0F83C3871C738CE6672666C9B24925B4B5AD4AD56AAAAAAAAAB55AB52969692DB6C9B266CCCC66318C71C7870F83E03FC001FFFFFE001FE03F0F87871E31C63198CCCCD99364934925A5A52B52A554AAAAAAAAB556AD4AD69696D24936C9B3266667339CE71C71E3C3E1F03F807FFE0000007FFC03F81F0787871E38C739CCE666666CD9B6492492DA5AD6B52B5";
defparam ram_block1a99.mem_init1 = "4AAB555555556AA956AD4A52D2D25B6DB649B3666CCCC667318E71C71E3C3C3E0F81FE00FFFC000000FFFE00FE07E0F87878F1C71C6318C6673333266CD936492492DA5A5AD6B52B54AAD5555AAAB55556AA55AB5A94B5A5B496DB6DB26C9B3266666663319CE31C63871E3C3C3E0F81F807FC003FFFFFFFFFFC001FF01FC1F83C1E1E3C78E38E31CE7319CCCCCCCCCD99364D924DB6925B4B6B4B5AD4AD5AB55AAA55555555555556AA954AB52B5294A5A5A5A4B6DB6DB6C9364C9933366666633398CE739C638E38E1C387878783E0FC1FC07F801FFE000000FFF8000007FFC00FF01F80F83E0F8787878F1E38F1CE38C739CE73399CCCCE664CCCD993264D";
defparam ram_block1a99.mem_init0 = "936C936DB6DB492DA5B4B4A5AD294AD4AD4A956AB556AAB55555AAAAAAAA955554AAAD54AA55AA54AD4AD6B5AD29694B69692DA492DB6DB6C926D936C99366CC99B33326666667333399CCE6339CE739C638C71C73871C70E3C78F0E1E1E1F0F0783E0F81F03F03F81FE03FC01FF800FFF80007FFFFF0000000000000001FFFFFC0001FFF000FFC00FF807F80FE03F81F81F81F03E0F83E0F0783C1E1E1F0F1E1E1E3C3870E1C78F1C78E38F1C71C71C738E38C718E31CE31CE718C639CE7318C67398C67319CC663319CCC66333999CCCC66673333399999998CCCCCCCCCCCCCCCCCCCCCCCD99999999B333333666666CCCCD9999B33326666CCCC9999B3336";

cyclonev_ram_block ram_block1a123(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a123_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a123.clk0_core_clock_enable = "ena0";
defparam ram_block1a123.clk0_input_clock_enable = "ena0";
defparam ram_block1a123.clk0_output_clock_enable = "ena0";
defparam ram_block1a123.data_interleave_offset_in_bits = 1;
defparam ram_block1a123.data_interleave_width_in_bits = 1;
defparam ram_block1a123.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a123.init_file_layout = "port_a";
defparam ram_block1a123.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a123.operation_mode = "rom";
defparam ram_block1a123.port_a_address_clear = "none";
defparam ram_block1a123.port_a_address_width = 13;
defparam ram_block1a123.port_a_data_out_clear = "none";
defparam ram_block1a123.port_a_data_out_clock = "clock0";
defparam ram_block1a123.port_a_data_width = 1;
defparam ram_block1a123.port_a_first_address = 40960;
defparam ram_block1a123.port_a_first_bit_number = 3;
defparam ram_block1a123.port_a_last_address = 49151;
defparam ram_block1a123.port_a_logical_ram_depth = 65536;
defparam ram_block1a123.port_a_logical_ram_width = 24;
defparam ram_block1a123.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a123.ram_block_type = "auto";
defparam ram_block1a123.mem_init3 = "000FE0F1C73999936DA5AD4AAAAAB56B496C993198E38783FE0001FF07871C673264DB4B5A9555554A94B6DB2666739E3C1F80000007E1E1C633333649696A55555552B4B4936666631C3C3F8000000FC1E38E733326DB694A9555554A9696DB3666338E1E0FE000003F83C38C633364DA4B5AB555556AD696D93666318E1E0FC000001FC1E38E733336496D6A556AAD54A52DB64CCCCE71E1E03FFFFFF80F0F1CE66664DB694A552AAB55A96924993318C71E0F800FFC00FC3C39C66664DB6D2952AAAAAB5296D36CCCCC638F0F807FFFF00F878E398CC992496B5AA9552AB5292DB26666738F0F03FF003FF83E1C719CCC9B25B4AD5AAAAA95296924D9999C";
defparam ram_block1a123.mem_init2 = "E38783F800000FE0F0E39CCCCD924B4A54AAAAA95296924D9999CE38783F8000007F078E38CE64C9B69695AAB54AA95AD2493666731C70F81FFC07FF81E1E39CC66CD92DA52B5555554AD69249B33339C71F0FE0000007F078E38CC64C9B69695AA9552AB5296DB66CCC671C783E007FFC00F83C71CC6664DB6D2D4AA5555AA5696936CCCCC638F0F80FFFFFF80F870E73999B26DA5AD4AAAAAAB5296924D9999CE38F07E007FE003F0F0E398CCC9B25B4A54AAAAAAD5AD25B26CCCC638E1F07FC0003FE07871C6333326DB4B4AD552A555A9496DB26666318F0F07F800003FC1E1C718CCCC9B6D2D2B554A9556A52DA6D9B3398C70F0FC00FFF801F878718C6";
defparam ram_block1a123.mem_init1 = "666C924B5AD52AAAAD529496D93666739C78781FF8001FF03E1C718CCCCD924B4B52AAD56AAD4A5B6DB3667318E1C1F01FFFFFE03E0E1C63199B36CB696A552AAA954AD2DA4D933319C71E1F01FFFFFFC07C3C71CE6666C924B4A54AAAAAAD5AD6D24D9B3398C70F0F807FFFFF80F83C71CC6666C9B496B52A95552AB52D2DB64CD8CC638F0F83FF0001FF03E1E39C6666649B696B5AA95556AB5296DB6C99998C71C7C3F001FFE003F078E38C66666C925B5AD5AAAAAA95294B6DB26666631C78781FC000007F81E1E39CE6666C9B69694AB555555AA52D2DB64CCCCC638E1E07E00000007F07871C63399326DB696B52AAD54AA95AD2DA6D9B3319C63C783F";
defparam ram_block1a123.mem_init0 = "003FFFC00FC1E3C6398CCD9B24B694AD52AAAAD56A52DA4DB3666338C78F07E01FFFFF807E0F1C718CE64CDB25B4A52AD555556A94A5B49B664CC6738E1E1F80FFFFFFF80F83C71C63333364DB496B52A955556AB52969249B3263318E38783F00FFFFFC01F83C78E739999936CB696B52A955556AB52969249B3666339C71E1F03FE00000FF81F0F1C719CCCCD936DA5A52A555595552A5296D26D9B33318C71C3C1F807FFFFFE01F07871C7399999B24925A5A952AAAAAAB56A5A5B6DB266666318E1C3C0FC001FF8007F07C38718C666664D924B4B5AB552AAAB552B5AD24924C99998C638E1E1F01FFE000FFF03F0F0E38C6733366C9249694AD56AAAAAA";

cyclonev_ram_block ram_block1a147(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a147_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a147.clk0_core_clock_enable = "ena0";
defparam ram_block1a147.clk0_input_clock_enable = "ena0";
defparam ram_block1a147.clk0_output_clock_enable = "ena0";
defparam ram_block1a147.data_interleave_offset_in_bits = 1;
defparam ram_block1a147.data_interleave_width_in_bits = 1;
defparam ram_block1a147.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a147.init_file_layout = "port_a";
defparam ram_block1a147.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a147.operation_mode = "rom";
defparam ram_block1a147.port_a_address_clear = "none";
defparam ram_block1a147.port_a_address_width = 13;
defparam ram_block1a147.port_a_data_out_clear = "none";
defparam ram_block1a147.port_a_data_out_clock = "clock0";
defparam ram_block1a147.port_a_data_width = 1;
defparam ram_block1a147.port_a_first_address = 49152;
defparam ram_block1a147.port_a_first_bit_number = 3;
defparam ram_block1a147.port_a_last_address = 57343;
defparam ram_block1a147.port_a_logical_ram_depth = 65536;
defparam ram_block1a147.port_a_logical_ram_width = 24;
defparam ram_block1a147.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a147.ram_block_type = "auto";
defparam ram_block1a147.mem_init3 = "AAAAAAD56A52D24926CD999CC638E1E1F81FFE000FFF01F0F0E38C6333326492496B5A955AAAA955AB5A5A49364CCCCC631C387C1FC003FF0007E07870E318CCCCC9B6DB4B4AD5AAAAAAA952B4B49249B333339C71C3C1F00FFFFFFC03F07871C631999B36C96D294A955535554A94B4B6D936666731C71E1F03FE00000FF81F0F1C7398CCD9B2492D295AAD55552A95AD2DA6D9333339CE3C783F007FFFFE01F83C38E3198C99B2492D295AAD55552A95AD25B64D99998C71C783E03FFFFFFE03F0F0E39CC664CDB25B4A52AD555556A94A5B49B664CE631C71E0FC03FFFFF00FC1E3C6398CCD9B64B694AD56AAAA956A52DA49B3666338C78F07E007FFF801";
defparam ram_block1a147.mem_init2 = "F83C78C73199B36CB696B52AA556AA95AD2DB6C993398C71C3C1FC0000000FC0F0E38C666664DB69694AB555555AA52D2DB26CCCCE738F0F03FC000007F03C3C718CCCCC9B6DA52952AAAAAB56B5B4926CCCCC638E3C1F800FFF001F87C71C6333326DB6D295AAD5552AB5AD2DB24CCCCC738F0F81FF0001FF83E1E38C663664DB69695AA95552A95AD25B26CCCC671C783E03FFFFFC03E1E1C63399B36496D6B56AAAAAA54A5A4926CCCCE71C787C07FFFFFF01F0F1C731999364B696A552AAA954AD2DA6D9B3318C70E0F80FFFFFF01F070E319CCD9B6DB4A56AAD56AA95A5A4936666631C70F81FF0003FF03C3C739CCCD936D252956AAAA956B5A4926CCC";
defparam ram_block1a147.mem_init1 = "C631C3C3F003FFE007E1E1C63399B36CB694AD552A555A9696DB2666631C70F07F800003FC1E1E318CCCC9B6D252B554A9556A5A5B6C99998C71C3C0FF80007FC1F0E38C6666C9B496B56AAAAAA54A5B49B2666338E1E1F800FFC00FC1E38E733336492D295AAAAAAA56B4B6C9B3339CE1C3E03FFFFFE03E1E38C66666D92D2D4AB5554AA5696DB64CCC671C783E007FFC00F83C71CC666CDB6D295AA9552AB52D2DB264C6638E3C1FC000000FE1F1C739999B2492D6A5555555A94B69366CC6738F0F03FFC07FF03E1C719CCCD92496B52AA55AAB52D2DB264CE638E3C1FC000003F83C38E733336492D2952AAAAA54A5A4936666738E1E0FE000003F83C38E";
defparam ram_block1a147.mem_init0 = "733336492D2952AAAAB56A5B49B266731C70F83FF801FF81E1E39CCCCC9B69295AA9552AB5AD2493266338E3C3E01FFFFC03E1E38C66666D96D295AAAAAA95296DB64CCCC738787E007FE003E0F1C6319932492D2B55AAA954A52DB64CCCCE71E1E03FFFFFF80F0F1CE66664DB694A556AAD54AD6D24D9999CE38F07F0000007E0F0E318CCD936D2D6AD55555AB5A4B64D998C638783F800000FE0F0E398CCD9B6D2D2A5555552A52DB6C9999CE38F07E0000003F878718CCCCD925A5A95555554AD2D24D99998C70F0FC0000003F078F39CCCC9B6DA52A5555552B5A5B64C99CC71C3C1FF0000FF83C38E3319326D25AD5AAAAAA56B4B6D933339C71E0FE000";

cyclonev_ram_block ram_block1a171(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a171_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a171.clk0_core_clock_enable = "ena0";
defparam ram_block1a171.clk0_input_clock_enable = "ena0";
defparam ram_block1a171.clk0_output_clock_enable = "ena0";
defparam ram_block1a171.data_interleave_offset_in_bits = 1;
defparam ram_block1a171.data_interleave_width_in_bits = 1;
defparam ram_block1a171.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a171.init_file_layout = "port_a";
defparam ram_block1a171.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a171.operation_mode = "rom";
defparam ram_block1a171.port_a_address_clear = "none";
defparam ram_block1a171.port_a_address_width = 13;
defparam ram_block1a171.port_a_data_out_clear = "none";
defparam ram_block1a171.port_a_data_out_clock = "clock0";
defparam ram_block1a171.port_a_data_width = 1;
defparam ram_block1a171.port_a_first_address = 57344;
defparam ram_block1a171.port_a_first_bit_number = 3;
defparam ram_block1a171.port_a_last_address = 65535;
defparam ram_block1a171.port_a_logical_ram_depth = 65536;
defparam ram_block1a171.port_a_logical_ram_width = 24;
defparam ram_block1a171.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a171.ram_block_type = "auto";
defparam ram_block1a171.mem_init3 = "D999B33326666CCCC9999B333366666CCCCCD999999B333333336666666666666666666666663333333399999CCCC6667333998CC6673198CC67319CC6339CC6319CE738C631CE718E718E31C638E39C71C71C71E38E3C71E3C70E1C3878F0F0F1E1F0F0F0783C1E0F83E0F81F03F03F03F80FE03FC03FE007FE001FFF00007FFFFF0000000000000001FFFFFC0003FFE003FF007F80FF03F81F81F03E0F83C1E1F0F0F0E1E3C78E1C71C39C71C638C739CE7398CE67339999CCCCCCC9999B3266CD9326D936C926DB6DB6924B692D2DA52D296B5AD6A56A54AB54AA556AAA555552AAAAAAAB55555AAAD55AAD52A56A56A5296B4A5A5B4B6925B6DB6D926D93";
defparam ram_block1a171.mem_init2 = "64C993366664CCE66673399CE739C638E71E38F1E3C3C3C3E0F83E03F01FE007FFC000003FFE000000FFF003FC07F07E0F83C3C3C3870E38E38C739CE633998CCCCCD9993264D926DB6DB6DA4B4B4B4A5295A95AA552AAD5555555555554AAB55AB56A56B5A5ADA5B492DB649364D9336666666667319CE718E38E3C78F0F0783F07F01FF0007FFFFFFFFFF8007FC03F03E0F87878F1C38C718E73198CCCCCCC99B26C9B6DB6D25B4B5A52B5AB54AAD5555AAAB55556AA55A95AD6B4B4B6924924D9366CC99999CCC6318C71C71E3C3C3E0FC0FE00FFFE0000007FFE00FF03E0F87878F1C71CE319CCC6666CCD9B24DB6DB4969694A56AD52AAD55555555AAA5";
defparam ram_block1a171.mem_init1 = "5A95AD6B4B6924924DB366CCCCCCE6739C638F1C3C3C1F03F807FFC000000FFFC03F81F0F878F1C71CE7399CCCCC99B26D92496D2D2D6A56AD55AAAAAAAAA554A95A94B4B4925924D933666663318C718F1C3C3E1F80FF000FFFFFF0007F80F83E1C3C71C6318CC6666CC9B26DB692D2D295AB55AAAAAAAAAAD56A56B5A5B49249B26CCC9CCCE639C71C38783E07E007FFFFFFFF801F81F07870E38C7399CCCCD9B36C925B4B4A52B54AAB55555AAAD5AB5A52DA4926D93366663318E71C38787C1FC03FFFFFFFFF807F07C3C38E38E73199999326D925B494B52B54AAAAAAAAA956AD6B4B69249B264CCCC6631C71C787C1F00FFE000003FF80FC1E1E3C738C";
defparam ram_block1a171.mem_init0 = "67333366C9B6DB4B4A52A552AAAAAAA552A529692DB6C9B33663318C71C70F07C0FF800000000FF03E0F0E38E318CCCCCC9B24925A5AD6AD54AAAAAA556AD6B4B6924D9326667318E71E3C1E07F000FFFF8007F03E1E3C738C6633266C9B6DA5A52952AB555552AB56A5A5A4926C99B3198C638E1E1E07F001FFFF800FE07C3871C7399CCD9936492DA5295AAD5555552A95AD692DB64D993399CE71C3C3C1FC01FFFFFE00FE0F0F1E31CE666664D9249696B52AD5555554AB529696DB6CD999998C71C70F07E01FFFFFFFE03F07870E318CC66CC9B6DB4B4AD4AA95555AA95294B6926D9B33319CE38F0F07E01FFFFFFC03F07878E39CC6664C9B6DA4A52B54";

cyclonev_ram_block ram_block1a51(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a51_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a51.clk0_core_clock_enable = "ena0";
defparam ram_block1a51.clk0_input_clock_enable = "ena0";
defparam ram_block1a51.clk0_output_clock_enable = "ena0";
defparam ram_block1a51.data_interleave_offset_in_bits = 1;
defparam ram_block1a51.data_interleave_width_in_bits = 1;
defparam ram_block1a51.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a51.init_file_layout = "port_a";
defparam ram_block1a51.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a51.operation_mode = "rom";
defparam ram_block1a51.port_a_address_clear = "none";
defparam ram_block1a51.port_a_address_width = 13;
defparam ram_block1a51.port_a_data_out_clear = "none";
defparam ram_block1a51.port_a_data_out_clock = "clock0";
defparam ram_block1a51.port_a_data_width = 1;
defparam ram_block1a51.port_a_first_address = 16384;
defparam ram_block1a51.port_a_first_bit_number = 3;
defparam ram_block1a51.port_a_last_address = 24575;
defparam ram_block1a51.port_a_logical_ram_depth = 65536;
defparam ram_block1a51.port_a_logical_ram_width = 24;
defparam ram_block1a51.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a51.ram_block_type = "auto";
defparam ram_block1a51.mem_init3 = "5555554AB5AD2DA4DB36666739C71E3E0FC007FFFE007E0F870E718CCCCC9B249696B52A955555AAD5A52DB6D932667318E38787C07FE0001FFC0F87871C63319B324DB496B5AB55555554A94A5B4936CCD8CC631C387C0FE0000000FE07878E38C66666C9B6D2D2952AA555AAA56B5B4924D99999CE71E3E1F807FFFFF803F0F0E38E6333366DB6D2D2B55AAAAAB54AD692DB64CCCCCE71C787C1FE000000FF03C3C71C6733366DB6D2D2B54AAAAA954A52D249366666739C38783F80000000FE0F871C631999B26DB4B4AD5AAAAAAB56A5A5B6C9B33398C71E1E07F8000007F81E1E38C6333364DB69695AA555554AB52D2DB6CD9998C638F0F03FE00001FF";
defparam ram_block1a51.mem_init2 = "03C3C718C6666C9B6D2D6A556AAAD54AD692DB264CCE639C3C3E07FFFFFFF81F0F1C7198CD9B2492D2B56AAAAAAD5A969249B327339C70E0F80FFFFFFC07E1E38E33999324925A52A5555555AB5A5B6D93263318E3C3E0FFC0003FF07C3C738CCCCC9B6D2D2B54AAAAB54AD6D249B366339C70F0FC01FFFF807E0F1C719CCC992492D6B55AAAAB54AD2D249B333318E38783F8000000FE0F0E38CE666CDB6D2D6AD5555552B5ADB4D9333338C78F07F00000007F0F8E38C6666CDB69294AB55555AA5292DB66CCCC638E1E0FE0000007F07871C6733364DB4B4AD54AAAD54A52DB6D9B3398E78F0FC01FFFF007C1E38E7333364925A52AD55554AB5A5B6D9333";
defparam ram_block1a51.mem_init1 = "318E387C1FF00007FC1F0E38CE666CDB69695AA9554AA56B4924D99998C70E1F80FFFFFE01F0F1C6339B324D25AD6AA5552AB5AD24926666631C383E01FFFFE01F0F1E739999B249694AD5555552B5A5B6C99998C71C3C0FF8000FF81E1C31CCCCC9B6DA52B555A5552B5B4926CCCCE71C3C1F8000000FE0F1C719CC9936DA5A956AAAAD529496C9B33318C38781FE0000FF03C38E31999B2492D2B55AAAB55A96924993339CE3C3E07FFFFFF81F0E18E63366C92D2D5AAAAAAAD4A4B6D9B3339C71E0F801FFE007E1E38E733326CB696A552AAB55A96924993339CE3C3E07FFFFFE03E1C71CCE4CDB6DA52A5555552A52DB6D99399C61C3E03FFFFFE03E1C31";
defparam ram_block1a51.mem_init0 = "CCE4CDB6DA52A555555AB5A5B6C9999CE38F0FC01FFF803F0F1C7319932492D2B55AAAB55AD2DA6C9998C638783FC00001FC0F1E719CCD936D2D2B5555554A9696D9333339C70F83FE0007FC0F0E38C6664DB6DAD6AB5554AA52D2493266338E3C1F800FE003F078E398CC99249695AA5554AA5696DB264C6738F0F01FFFFFFC0F871C633336492D2D5AAAAAAD5A5A493666631C78780FFFFFF80F871C6333364925AD4AAAAAA952D2DB26666738F1F03FFC0FFE07C38E3399B36DB4A52AA552AA5296DB66CCE638E1F07FF80FFE07C78E7333326DA5AD4AAAAAA95AD2493266739C387E03FFFFC07E1C39CE664C925A5AB5555552B5A4924CCCCE31E1E03FFF";

cyclonev_ram_block ram_block1a75(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a75_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a75.clk0_core_clock_enable = "ena0";
defparam ram_block1a75.clk0_input_clock_enable = "ena0";
defparam ram_block1a75.clk0_output_clock_enable = "ena0";
defparam ram_block1a75.data_interleave_offset_in_bits = 1;
defparam ram_block1a75.data_interleave_width_in_bits = 1;
defparam ram_block1a75.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a75.init_file_layout = "port_a";
defparam ram_block1a75.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a75.operation_mode = "rom";
defparam ram_block1a75.port_a_address_clear = "none";
defparam ram_block1a75.port_a_address_width = 13;
defparam ram_block1a75.port_a_data_out_clear = "none";
defparam ram_block1a75.port_a_data_out_clock = "clock0";
defparam ram_block1a75.port_a_data_width = 1;
defparam ram_block1a75.port_a_first_address = 24576;
defparam ram_block1a75.port_a_first_bit_number = 3;
defparam ram_block1a75.port_a_last_address = 32767;
defparam ram_block1a75.port_a_logical_ram_depth = 65536;
defparam ram_block1a75.port_a_logical_ram_width = 24;
defparam ram_block1a75.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a75.ram_block_type = "auto";
defparam ram_block1a75.mem_init3 = "6664CCCD999B333266664CCCD99999333336666664CCCCCCCD99999999999999999999999999998CCCCCCE66663333999CCCE6633399CCE63319CC67318CE7318C6318C6318E738C738C738E31C738E38E38E38E38F1C78E3C70E1C3878F0F1E1E1E1E1F0F0783C1F0F83F07C0F81F81F80FE03F807F803FF003FF8003FFFC00000FFFFFFFFFFFFFFFFFE000007FFF000FFE007FC03F807E03F03F07C0F87C1E0F0F0F0F0E1E3C70E3871C71C638E718C739CC63399CCE6673333333332666CC99B364D93649B64924924925B692D25A5A5AD296B5A94AD5A956A956AAD556AAAAD5555555554AAAA9554AAD56A952B52B5AD6B5A5A5A5A4B6D24924924DB24D";
defparam ram_block1a75.mem_init2 = "93264C999B3333331998CE6339CE31C638E3871E3C78787C3E0F81F81FC03FF000FFFFF0000003FFFFC003FE01FC0FC0F83C1E1E1C3871C71C718E7398CE6633333332664C9B26C926DB6D24B69696B4A52B52A54AA555AAAAAA55AAAAAA555AAD5AB5294A52D2D25B4924926D9364CD99B3333999CC6738C71C71C78F0F0F07C1F81FC01FFE000000000001FFE01FC07E0F8783878F1C71CE318C6733333333266C9B24936925B4B4B5AD6A56A955AAAA555554AAAB552AD4AD6B4A5B4B6DB6DB64D9B326666663318C638C70E3C787C3E07E03FE000FFFFFFFF0007F807E0F83C3C78E38E39CE7339999993364D92492496D2D6B5AD5AA554AAAAAAAAA9552";
defparam ram_block1a75.mem_init1 = "AD4AD6B4B4B6D249B64D9B333333398CE31C71C3C783C0F80FF000FFFFFFFE001FE03E0F87878E38E39CE6733333266C9B6DB6D25A5294AD5AA95555555556AA54AD6B5A4B69249B66CD999998CC639C71C3C7C3E0FE03FFC0000001FFC03F03E1E1E38E38C633999999326C92492DA5AD6B56A95554AAD5556AB52B5A5A5B6DB6C9B326667339CE31C3878783F03FE0000000001FE03F0787871C718C673333366C9B6DB49694A56A9552AAAAAB556AD4A52D2DB6DB26CD99998CE738E3870F07C07F80007FC0003FC0FC3E3C78E318C6666664C936DB49694A56A95552AA5554AB5294B4B6DB6C993333339CE71C38787C0FE007FFFFFF003F83E0F1E38E71";
defparam ram_block1a75.mem_init0 = "9CCCCCD9B24924B6B4AD4AA555555552A95A96B6924926CC9999CC631C78F0F07E01FFFFFFFFF807E0F0F0E38C633199B326D92DB4B5AD5AAD5555552AB52B4B4B6DB64C99999CC638E3C3C1F01FFC00001FFC07C1E1E38E719CCCCD9B24924B4A52A556AAAAAB55AB5AD2DB6DB264CCCE631C71C3C1F01FF800001FF80F83C38718C67333264DB6DA5A52B54AAAAAAAB54AD6969249366CCCC6738E38787E07FC000000FF81F87871C63198CD9936DB6D296A55AAAAAAAA55A94B496C9366CCC6739C70F0F03F800000000FE07C3871C633999B364DA496B5A955AAAAA954A94B4B6DB26CCCCC671C71E1F03FC0000001FE07C3C71C6319999324924B4A56A9";

cyclonev_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 8191;
defparam ram_block1a3.port_a_logical_ram_depth = 65536;
defparam ram_block1a3.port_a_logical_ram_width = 24;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init3 = "2AD4A5A492499333318C71C787C0FF00000007F81F0F1C71CC66666C9B6DA5A52A552AAAAB552B5AD24B64D9B33398C71C387C0FE000000003F81E1E1C739CC666CD926D25A52B54AAAAAAAB54AD296DB6D933663318C71C3C3F03FE0000007FC0FC3C38E39CC6666CD92492D2D6A55AAAAAAAA55A94B4B6DB64C9999CC631C38783E03FF000003FF01F07871C718CE6664C9B6DB696B5AB55AAAAAAD54A94A5A49249B36666731CE38F0F07C07FF000007FF01F07878E38C673333264DB6DA5A5A95AA95555556AB56B5A5B6936C99B33198C638E1E1E0FC03FFFFFFFFF00FC1E1E3C718C67333266C92492DAD2B52A955555554AA56A5ADA49249B36666673";
defparam ram_block1a3.mem_init2 = "1CE38F1E0F83F801FFFFFFC00FE07C3C3871CE73999999326DB6DA5A5295AA5554AA95552AD4A52D25B6D9264CCCCCC6318E3C78F87E07F80007FC0003FC07C1E1C38E39CE63333366C9B6DB69694A56AD55AAAAAA9552AD4A52D25B6DB26CD99999CC631C71C3C3C1F80FF0000000000FF81F83C3C38718E7399CCCC99B26DB6DB4B4B5A95AAD5556AA55552AD5AD6B4B6924926C9933333398C638E38F0F0F81F807FF00000007FF80FE0F87C7871C738C6633333366CDB2492DA4B5AD6A54AAD5555555552AB56A5294B496DB6DB26CC999999CCE738E38E3C3C3E0F80FF000FFFFFFFE001FE03E0783C7871C718E6339999999B364DB2496DA5A5AD6A56A";
defparam ram_block1a3.mem_init1 = "9552AAAAAAAAA554AB56B5AD696D249249364D9933333399CE738E38E3C78783E0FC03FC001FFFFFFFE000FF80FC0F87C3C78E1C638C63198CCCCCC99B364DB6DB6DA5B4A5AD6A56A955AAAA555554AAAB552AD4AD6B5A5A5B492D9249B26CC999999999CC6318E71C71E3C383C3E0FC07F00FFF000000000000FFF007F03F07C1E1E1E3C71C71C639CC673339999B33664D936C924925B4969694A5295AB56AB554AAAAAB54AAAAAB554AA54A95A94A5AD2D2DA496DB6C926C9B264CC99999998CCE6339CE31C71C71C3870F0F0783E07E07F00FF8007FFFF8000001FFFFE001FF807F03F03E0F87C3C3C78F1C38E38C718E7398CE63331999999B33264C993";
defparam ram_block1a3.mem_init0 = "649B6492492496DA4B4B4B4B5AD6B5A95A952AD56AA5552AAAA55555555556AAAAD556AAD52AD52B56A52B5AD296B4B4B49692DB4924924924DB24D9364D9B3266CCC9999999999CCCE673398C6739C631CE38C71C71C38E1C78F0E1E1E1E1E0F07C3E07C1F81F80FC03F807FC00FFE001FFFC00000FFFFFFFFFFFFFFFFFE000007FFF8003FF801FF803FC03F80FE03F03F03E07C1F83E1F0783C1E1F0F0F0F0F1E1E3C3870E1C78E3C71E38E38E38E38E39C718E39C639C639CE318C6318C6319CE6319CC673198CE6733998CCE6673339998CCCCE66666633333333333333333333333333333666666664CCCCCD999993333366664CCCC9999B33366664CCC";

cyclonev_ram_block ram_block1a27(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.clk0_output_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "rom";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "clock0";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 8192;
defparam ram_block1a27.port_a_first_bit_number = 3;
defparam ram_block1a27.port_a_last_address = 16383;
defparam ram_block1a27.port_a_logical_ram_depth = 65536;
defparam ram_block1a27.port_a_logical_ram_width = 24;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init3 = "FFF80F0F18E66664924B5A9555555AB4B49264CCE73870FC07FFFF80FC38739CCC992496B52AAAAAA56B4B6C99999CE3C7C0FFE03FFC1F0E38CE66CDB6D294AA954AA94A5B6D9B3398E387C0FFE07FF81F1E39CCCCC9B696952AAAAAA56B4924D9998C71C3E03FFFFFE03C3C718CCCD924B4B56AAAAAB5696924D9998C71C3E07FFFFFF01E1E39CC64C9B6D2D4AA5554AB52D2493266338E3C1F800FE003F078E398CC99249694AA5555AAD6B6DB64CCC638E1E07FC000FF83E1C739999936D2D2A5555555A9696D9366731CF1E07F000007F83C38C633326CB696B55AAAB55A96924993319C71E1F803FFF007E1E38E733326DB4B5AB555554A94B6DB664E67";
defparam ram_block1a27.mem_init2 = "1870F80FFFFFF80F870C7339336DB694A9555554A94B6DB664E671C70F80FFFFFFC0F878E7399932492D2B55AAA954AD2DA6C9999CE38F0FC00FFF003E0F1C73999B36DA4A56AAAAAAB5696926CD98CE30E1F03FFFFFFC0F878E7399932492D2B55AAAB55A969249B33318E38781FE0000FF03C38631999B26D252956AAAAD52B4B6D9326731C71E0FE0000003F07871CE6666C925B5A9554B555A94B6DB2666671870F03FE0003FE07871C6333326DB4B5A95555556A52D249B33339CF1E1F00FFFFF00F838718CCCCC92496B5AA9554AAD6B496499B398C71E1F00FFFFFE03F0E1C63333364925AD4AA5552AB52D2DB66CCCE638E1F07FC0001FF07C38E319";
defparam ram_block1a27.mem_init1 = "99936DB4B5AA555556A94B4924D9999CE38F07C01FFFF007E1E3CE3399B36DB694A556AAA556A5A5B64D999CC71C3C1FC000000FE0F0E38C6666CDB69294AB55555AA5292DB66CCCC638E3E1FC0000001FC1E3C6399999365B6B5A95555556AD696DB66CCCE638E1E0FE0000003F83C38E319999B249696A55AAAAB55AD692493266731C71E0FC03FFFF007E1E1C7398CD9B2496D6A55AAAAA55A9696DB26666639C787C1FF80007FE0F878E3198C9936DB4B5AB5555554A94B49249933398E38F0FC07FFFFFE03E0E1C7399C99B2492D2B56AAAAAAD5A969249B366331C71E1F03FFFFFFFC0F878738CE664C9B692D6A556AAAD54AD696DB26CCCC631C78781";
defparam ram_block1a27.mem_init0 = "FF00000FF81E1E38C6333366DB69695AA555554AB52D2DB64D9998C638F0F03FC000003FC0F0F1C633999B26DB4B4AD5AAAAAAB56A5A5B6C9B33318C71C3E0FE00000003F83C38739CCCCCD9249694A552AAAAA55A9696DB6CD999CC71C78781FE000000FF07C3C71CE666664DB692D6A55AAAAAB55A9696DB6CD9998CE38E1E1F803FFFFFC03F0F8F1CE73333364925B5AD4AAB554AA9529696DB26CCCCC638E3C3C0FE0000000FE07C38718C663666D925B4A52A55555555AB5AD25B6499B3198C71C3C3E07FF0000FFC07C3C38E319CCC9936DB694B56AB555552A95AD2D249B26666631CE1C3E0FC00FFFFC007E0F8F1C739CCCCD9B64B696B5AA5555555";

cyclonev_ram_block ram_block1a100(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a100_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a100.clk0_core_clock_enable = "ena0";
defparam ram_block1a100.clk0_input_clock_enable = "ena0";
defparam ram_block1a100.clk0_output_clock_enable = "ena0";
defparam ram_block1a100.data_interleave_offset_in_bits = 1;
defparam ram_block1a100.data_interleave_width_in_bits = 1;
defparam ram_block1a100.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a100.init_file_layout = "port_a";
defparam ram_block1a100.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a100.operation_mode = "rom";
defparam ram_block1a100.port_a_address_clear = "none";
defparam ram_block1a100.port_a_address_width = 13;
defparam ram_block1a100.port_a_data_out_clear = "none";
defparam ram_block1a100.port_a_data_out_clock = "clock0";
defparam ram_block1a100.port_a_data_width = 1;
defparam ram_block1a100.port_a_first_address = 32768;
defparam ram_block1a100.port_a_first_bit_number = 4;
defparam ram_block1a100.port_a_last_address = 40959;
defparam ram_block1a100.port_a_logical_ram_depth = 65536;
defparam ram_block1a100.port_a_logical_ram_width = 24;
defparam ram_block1a100.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a100.ram_block_type = "auto";
defparam ram_block1a100.mem_init3 = "66318C738E3C78F0F87C0FC03FE0007FFFFFF0003FE01F81F0F87870E38E39CE73198CCCC999326C936DB692DA52D6B5AB56AB555AAAAAAAA5556AB56A56B5A5A5A4B6DB649B26CC99999998CE631CE38E3870F0F0F81F01FE00FFFF000000FFFF007F80FC1F0F870F1C38E71CE73198CCCCCCD99364D924924B692D296B52B56AD55AAAA95555AAAA955AA54AD6B5A52DA4B6DB6D926C99332666663319CE738C71C38F0E1F0F83E07F00FFE00003FFFE00003FF007F03E0F83C3C78F1C71C639CE633399999933264D926DB6DB692D2D2D6B5A95AB55AAB5555555555554AA954A95A94A52D692D24B6DB249B26CD993333333198CE739C638E3C70E1E1E0F";
defparam ram_block1a100.mem_init2 = "83E07F00FF8003FFFFFFFFFFE000FFC03F03F07C3E1E1C3871C71C639CE63319999999993364C936C924925B4969694B5A95A952AD54AAA95555555552AAA556A952A56B5AD29696D25B6DB6DB26D93264CCD99999CCC66318C639C71C71E3C78787C3E07C0FE03FE003FFFC000000003FFFC007FC07F03F07C1E1F1E1E3871C71C738C6339CCE6666666666CC99364DB249B6DA496D25A5AD294A52B52AD5AA9556AAAAB555554AAAAB555AAD52A54A56B5AD2969692DA4925924936C9B264C999333333333998CE7318E718E38E38F1C3C78787C3E0F81F81FC03FE003FFF80000000000003FFF800FF807F01F83F07C3E1E1E1E3C78E38E38E39C6318CE73";
defparam ram_block1a100.mem_init1 = "3998CCCCCCCCD99B3264D93649B6C92492DB692D25A5AD2D6B5AD4AD4A956A955AAB5555AAAAAAAAAAAAAB5554AAB552AD52A56A56B5AD6B4A5A5A4B496DA4924924936C9364D9B266CC99999333399998CC66339CE739C638E71C71C38F1C3C7878787C3E1F03E07C07E03FC03FF001FFF800003FFFFFFFFFFC00000FFFC007FC01FE03F81F81F03E0F07C3C3C3C3C3870E3C71C38E71C738E738C6339CC6733999CCCCCCCCCCCCCD99B3266C99364D936C936D924924925B6D25B49692D2D2D696B5A5294AD6A56A54A952AD52A955AAB5552AAAB555555555AAAD555555556AAAA5552AAD54AAD52AD52A54AD5A94AD6A5294A5AD29696B4B69696D25B496";
defparam ram_block1a100.mem_init0 = "DA4925B6DB6D924936D926C9364D9366C993264CD99B33266666CCCCCCCCE66667333198CC663398CE7318C631CE718C718E31C71CE38E38F1C71E38F1E3870F1E3C3C387878783C3C1E0F07C3E0F83E07C0F81F83F81F80FC07F00FE01FE00FF803FF001FFC003FFE0003FFFE00000FFFFFFF8000000000000000000000000003FFFFFFF000003FFFF80007FFE0007FF8007FF001FF801FF007FC01FE00FF01FE01FC07F01FC07F03F81F80FC0FC0FC0F81F83F07E0FC1F03E0F83E07C1F0F83E0F87C1F0F83C1E0F07C3C1E0F0787C3C3E1E0F0F0F87878787C3C3C3C3C3C3C3C3C3C3C3C3878787878F0F0F0E1E1E1C3C3C787870F0E1E1E3C3C787870F0E";

cyclonev_ram_block ram_block1a124(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a124_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a124.clk0_core_clock_enable = "ena0";
defparam ram_block1a124.clk0_input_clock_enable = "ena0";
defparam ram_block1a124.clk0_output_clock_enable = "ena0";
defparam ram_block1a124.data_interleave_offset_in_bits = 1;
defparam ram_block1a124.data_interleave_width_in_bits = 1;
defparam ram_block1a124.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a124.init_file_layout = "port_a";
defparam ram_block1a124.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a124.operation_mode = "rom";
defparam ram_block1a124.port_a_address_clear = "none";
defparam ram_block1a124.port_a_address_width = 13;
defparam ram_block1a124.port_a_data_out_clear = "none";
defparam ram_block1a124.port_a_data_out_clock = "clock0";
defparam ram_block1a124.port_a_data_width = 1;
defparam ram_block1a124.port_a_first_address = 40960;
defparam ram_block1a124.port_a_first_bit_number = 4;
defparam ram_block1a124.port_a_last_address = 49151;
defparam ram_block1a124.port_a_logical_ram_depth = 65536;
defparam ram_block1a124.port_a_logical_ram_width = 24;
defparam ram_block1a124.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a124.ram_block_type = "auto";
defparam ram_block1a124.mem_init3 = "00001FF03F07878F1C639CC666666CD924DA4B6B4A56AD56AAAAAAAA552A56B5A4B6926D932666667318C71C38787C1FC01FFFFFFFFFE01FC1F0F0F1C718E6333333366D92492D2D294A956AAAAAAAAA954AD4A5A5B4924D932666667318E71C38783C0FE00FFFFFFFFF803F83E0F0E3C638C6733333264DB24B6D2D6B5AB55AAAAAAAAA954AD4A5A5A49249B3664CCE6739CE3870F0F07E01FFC0000007FF00FC1E1E1C38E739CCE666CC9B24924B694A52B55AAAA556AAA956AD6B4B496DB64D9B3333339CE71C70F0F07C0FF0007FFFF0007F81F87C3871C718C66733666C9B6496D2D2D6A55AA955555552AB56A529692DB6D9366CCCCCE6318E38E1E1E0";
defparam ram_block1a124.mem_init2 = "FC07FC000000001FF01F83C3C38E38C63399999B364DB6DB4B4B5A952A9555555555AAD4AD6B496D24DB26CCD98CCE631C71C78783E07F001FFFFFFF801FE07C3E1C38E39CE7333333264DB6DB69696B52B55AAAAAAAAAA552B5296B692DB24D9332663339CE71C78F0F87E07FC0007FFC0007FC0FC3E1E3C71CE3399CCCC99324DB6DA5A5AD6A55AAA5555552AAD5AB5AD2D24B6C9366CCCCCCC6318E38E1E1E0FC0FF80007FE0000FF01F87C3C78E38C633999999B364936925A5AD6A54AAD55555554AAD5A94A5A5B4926D936664C666318E71C38787C1F00FF8000000003FE03F07C3C3871CE318CCC64CCD9364924B696B5AD5AA5555AAAD5552AD5AD6B";
defparam ram_block1a124.mem_init1 = "4B4924926C99B333319CE718E1C78783E07F801FFFFFFFF001FC0F83C3C38E38C73199CCD99B26C92496D2D6B5AB54AAB555554AAB54A94A52D25B6DB24C99B333198CE31C71E3C3E1F81FE001FFFFFFC003FC0FC1E1E1C71C739CC6666664C9B24924B696B5AD5AA5552AAAAAD552A95A96B4B492D924D9B326663339CE31C78F1F0F83F00FFC00000000FFE01F83E1E1E38718E73998CCCD99364DB6DA4B4B5AD4AD56AAAB554AAAA552B5294B4B4924926C9933333319CE738E3C78787C1F807FE0000000007FE01F83E1E1E38718E7398CCCCCC993649B6D25A5A5295AB552AAAAAAAAAA552A56B5AD25B4924DB264CC998CCE631CE38E1C3C1E07C07FC0";
defparam ram_block1a124.mem_init0 = "003FFFC0003FE03E0783C3871C718C63319999B326C9B6DB692D296A52A552AAB555552AAB55A95AD6B496924926C9B36666667318C638E3878F0783F01FE000FFFFFFF8007FC0FC1F0F0F1C38C718CE673333266C9B24924969296B5A952A9555AAAAA95552A952B5AD2D2DA4924DB264CD99998CC6318E38E3C787C3E07E01FFC0000000007FF00FC0F83C3C38F1C639CE63333B33366C9B24924B69694A52B56AB5552AAAAAB555AAD5A95AD2D2D24924936CD9B333333398C639C71C3878783E0FE03FF00001FF80000FFC07F07C1E1E1C38E38C7398CCE6666CC99364924925B4B4A5295AB54AAB555555555AAA55AB5294A5A5B4924924D93664CCCCCC";

cyclonev_ram_block ram_block1a148(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a148_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a148.clk0_core_clock_enable = "ena0";
defparam ram_block1a148.clk0_input_clock_enable = "ena0";
defparam ram_block1a148.clk0_output_clock_enable = "ena0";
defparam ram_block1a148.data_interleave_offset_in_bits = 1;
defparam ram_block1a148.data_interleave_width_in_bits = 1;
defparam ram_block1a148.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a148.init_file_layout = "port_a";
defparam ram_block1a148.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a148.operation_mode = "rom";
defparam ram_block1a148.port_a_address_clear = "none";
defparam ram_block1a148.port_a_address_width = 13;
defparam ram_block1a148.port_a_data_out_clear = "none";
defparam ram_block1a148.port_a_data_out_clock = "clock0";
defparam ram_block1a148.port_a_data_width = 1;
defparam ram_block1a148.port_a_first_address = 49152;
defparam ram_block1a148.port_a_first_bit_number = 4;
defparam ram_block1a148.port_a_last_address = 57343;
defparam ram_block1a148.port_a_logical_ram_depth = 65536;
defparam ram_block1a148.port_a_logical_ram_width = 24;
defparam ram_block1a148.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a148.ram_block_type = "auto";
defparam ram_block1a148.mem_init3 = "6666664CD9364924925B4B4A5295AB54AAB555555555AAA55AB5294A5A5B4924924D93266CCCCE66339C638E3870F0F07C1FC07FE00003FF00001FF80FE0F83C3C3871C738C6339999999B366D924924969696B52B56AB555AAAAAA9555AAD5A94A52D2DA49249B26CD999B9998CE738C71E3878783E07E01FFC0000000007FF00FC0F87C3C78E38E318C6633333664C9B64924B69696B5A952A95552AAAAB5552A952B5AD292D249249B26CC99999CCE631C63871E1E1F07E07FC003FFFFFFE000FF01F83C1E3C38E38C6319CCCCCCD9B26C92492D25AD6B52B55AAA955555AAA954A94AD29692DB6DB26C99B3333198C631C71C38783C0F80FF80007FFF800";
defparam ram_block1a148.mem_init2 = "07FC07C0F07870E38E718CE66332664C9B64925B496B5AD4A954AAAAAAAAAA955AB5294B4B496DB24D932666666339CE31C38F0F0F83F00FFC000000000FFC03F07C3C3C78E39CE731999999326C924925A5A5295A954AAAA555AAAAD56A56B5A5A4B6DB64D93366663339CE31C38F0F0F83F00FFE000000007FE01F83E1F1E3C718E73998CCC99B364936925A5AD2B52A9556AAAAA9554AB56B5AD2DA49249B264CCCCCC6739C71C70F0F07E07F8007FFFFFF000FF03F0F878F1C718E6331999B32649B6DB49694A52A55AAA555555AAA55AB5AD696D24926C9B336673319C638E3878783E07F001FFFFFFFF003FC0F83C3C70E31CE7319999B326C924925A5";
defparam ram_block1a148.mem_init1 = "AD6B56A95556AAB5554AB56B5AD2DA4924D936664C666318E71C38787C1F80FF8000000003FE01F07C3C3871CE318CCC64CCD936C925B4B4A52B56AA555555556AA54AD6B4B492D924D9B33333398C638E3C787C3F01FE0000FFC0003FE07E0F0F0E38E318C6666666CD926DA49696B5AB56AA9555554AAB54AD6B4B4B6DB64993266673398E71C78F0F87E07FC0007FFC0007FC0FC3E1E3C71CE73998CC9993649B692DAD295A954AAAAAAAAAB55A95AD2D2DB6DB64C9999999CE738E3870F87C0FF003FFFFFFF001FC0F83C3C71C718CE6633666C9B6496D25AD6A56AB5555555552A952B5A5A5B6DB64D9B3333398C638E3878783F01FF0000000007FC07E";
defparam ram_block1a148.mem_init0 = "0F0F0E38E318CE66666CD936DB692D294AD5AA955555552AB54AD69696D24DB26CCD99CCC631C71C387C3F03FC001FFFFC001FE07C1E1E1C71CE73999999B364DB6D25A5AD6AD52AAAD54AAAB55A94A52DA49249B266CCCE6739CE3870F0F07E01FFC0000007FF00FC1E1E1C38E739CCE664CD9B24924B4B4A56A552AAAAAAAAB55AB5AD696DA49B64C999999CC638C78E1E0F83F803FFFFFFFFE00FE0783C3871CE319CCCCCC99364925B4B4A56A552AAAAAAAAAD52A529696924936CD9999998CE31C71E1E1F07F00FFFFFFFFFF007F07C3C3871C6319CCCCCC9936C92DA4B5AD4A954AAAAAAAAD56AD4A5ADA4B649366CCCCCC6738C71E3C3C1F81FF00000";

cyclonev_ram_block ram_block1a172(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a172_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a172.clk0_core_clock_enable = "ena0";
defparam ram_block1a172.clk0_input_clock_enable = "ena0";
defparam ram_block1a172.clk0_output_clock_enable = "ena0";
defparam ram_block1a172.data_interleave_offset_in_bits = 1;
defparam ram_block1a172.data_interleave_width_in_bits = 1;
defparam ram_block1a172.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a172.init_file_layout = "port_a";
defparam ram_block1a172.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a172.operation_mode = "rom";
defparam ram_block1a172.port_a_address_clear = "none";
defparam ram_block1a172.port_a_address_width = 13;
defparam ram_block1a172.port_a_data_out_clear = "none";
defparam ram_block1a172.port_a_data_out_clock = "clock0";
defparam ram_block1a172.port_a_data_width = 1;
defparam ram_block1a172.port_a_first_address = 57344;
defparam ram_block1a172.port_a_first_bit_number = 4;
defparam ram_block1a172.port_a_last_address = 65535;
defparam ram_block1a172.port_a_logical_ram_depth = 65536;
defparam ram_block1a172.port_a_logical_ram_width = 24;
defparam ram_block1a172.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a172.ram_block_type = "auto";
defparam ram_block1a172.mem_init3 = "E1E1C3C3C7878F0F0E1E1C3C3C787870F0F0E1E1E1E3C3C3C3C3878787878787878787878787C3C3C3C3E1E1E0F0F8787C3C1E0F0787C1E0F0783E1F07C3E0F83E1F07C0F83E0F81F07E0FC1F83F03E07E07E07E03F03F81FC07F01FC07F00FF01FE00FF007FC01FF003FF001FFC003FFC000FFFC0003FFFF800001FFFFFFF8000000000000000000000000003FFFFFFE00000FFFF8000FFF8007FF001FF803FE00FF00FE01FC07E03F03F83F03E07C0F83E0F87C1E0F078783C3C3C387878F1E1C38F1E38F1C71E38E38E71C718E31C631CE718C6319CE63398CC66331999CCCCCE66666666CCCCC999B33664C99326CD9364D926C936D924936DB6DB4924B6";
defparam ram_block1a172.mem_init2 = "D25B496D2D2DA5AD2D296B4A5294AD6A52B56A54A956A956AA556AA9554AAAAD555555556AAB555555555AAAA9555AAB552A956A952A54AD4AD6A5294B5AD2D6969692D25B496DB4924924936D926D9364D9326CC99B336666666666666733399CC67398C639CE39C71CE3871C78E1C38787878787C1E0F81F03F03F80FF007FC007FFE000007FFFFFFFFFF800003FFF001FF807F80FC07C0F81F0F87C3C3C3C7871E3871C71CE38C739CE7398CC663333399993333266CC9B364D926D924924924B6D25A4B4B4A5AD6B5AD4AD4A956A955AAA5555AAAAAAAAAAAAAB5555AAB552AD52A56A56B5AD696B4B49692DB6924926DB24D9364C99B336666666663339";
defparam ram_block1a172.mem_init1 = "9CE6318C738E38E38E3C78F0F0F0F87C1F83F01FC03FE003FFF80000000000003FFF800FF807F03F03E0F87C3C3C7871E38E38E31CE319CE633399999999933264C9B26D924934924B692D2D296B5AD4A54A956AB555AAAAA555555AAAAAD552AB56A95A94A5296B4B496D24B6DB249B64D93266CCCCCCCCCCE67398C639C71C71C38F0F1F0F07C1F81FC07FC007FFF8000000007FFF800FF80FE07C0F87C3C3C78F1C71C738C6318CC667333336664C9936C9B6DB6DB496D2D296B5AD4A952AD54AAA95555555552AAA556A952B52B5A52D2D25B4924926D9264D99333333333198CE738C71C71C3870F0F87C1F81F807FE000FFFFFFFFFFF8003FE01FC0F83";
defparam ram_block1a172.mem_init0 = "E0F0F0E1C78E38C739CE633199999993366C9B249B6DA49692D694A52B52A552AA5555555555555AAB55AB52B5AD6969692DB6DB6C9364C999333333998CE738C71C71E3C78783E0F81FC01FF80000FFFF80000FFE01FC0F83E1F0E1E3871C639CE73198CCCCC999326C936DB6DA4B694B5AD6A54AB552AAAB55552AAAB556AD5A95AD29692DA49249364D93366666663319CE71CE3871E1C3E1F07E03FC01FFFE000001FFFE00FF01F03E1E1E1C38E38E718CE63333333266C9B24DB6DA4B4B4B5AD4AD5AAD554AAAAAAAB555AAD5AB5AD694B692DB6D926C9933266663319CE738E38E1C3C3E1F03F00FF8001FFFFFFC000FF807E07C3E1E3C78E39C6318CC";

cyclonev_ram_block ram_block1a52(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a52_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a52.clk0_core_clock_enable = "ena0";
defparam ram_block1a52.clk0_input_clock_enable = "ena0";
defparam ram_block1a52.clk0_output_clock_enable = "ena0";
defparam ram_block1a52.data_interleave_offset_in_bits = 1;
defparam ram_block1a52.data_interleave_width_in_bits = 1;
defparam ram_block1a52.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a52.init_file_layout = "port_a";
defparam ram_block1a52.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a52.operation_mode = "rom";
defparam ram_block1a52.port_a_address_clear = "none";
defparam ram_block1a52.port_a_address_width = 13;
defparam ram_block1a52.port_a_data_out_clear = "none";
defparam ram_block1a52.port_a_data_out_clock = "clock0";
defparam ram_block1a52.port_a_data_width = 1;
defparam ram_block1a52.port_a_first_address = 16384;
defparam ram_block1a52.port_a_first_bit_number = 4;
defparam ram_block1a52.port_a_last_address = 24575;
defparam ram_block1a52.port_a_logical_ram_depth = 65536;
defparam ram_block1a52.port_a_logical_ram_width = 24;
defparam ram_block1a52.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a52.ram_block_type = "auto";
defparam ram_block1a52.mem_init3 = "9999999326C9B6C96DA4B4B5AD6A54AB556AAAAAAAAAD55AAD5AD4A5A5A5B6924DB26C99B3333399CC631C71C70E1E0F07E07F803FFFE0001FFFF007F81F83C1E3C38E38E739CC66666666CD936D925B696D694A56AD56AAB5555555AAAD52A56A52D2D25B6DB649B3666CCC666318C738E3C78787C1F01FE007FFFFFFFFFC00FF03F07C3C3871C71CE3399CCCCCD99364DB6DB6969694A56AD56AAB555555AAA956AD4AD29692DB6DB649932666667339CE31C70E1E1E0F83F807FF80000000FFF007E07C1E1E3C71C738CE6333333264C936DB6D25A52D6A54AB5552AAAAAD554AB56A529696D24924DB366CCCCCC6731CE38E3C78783E07F00FFFE00001FF";
defparam ram_block1a52.mem_init2 = "FC03F81F07878F1C71CE73998CCC999364DB6DB49694B52956AB55555555554AA54AD4B5A4B69249B66CD999999CC6718E3870E0F07C0FE007FFFFFFFFF801FC0FC3E1E3C71C639CC6666666CD936DB6DA4B5A52B56AB5556AAA95552A95295A5A5A49249B66CD99998CC631CE3870E1F07C0FF003FFFFFFFF800FE07E1F0F1E38E318C663333266C9B6492DA5A5AD4AD52AAD555555AAA55A95A52D25B6DB64D9B33333318C638C38F0F0F83F80FFF00000007FF00FC0F87870E38E318CC66666CC9B24924B69694AD4AB554AAAAAAD552AD4AD29692DB6D9264CD999CCC631C71C78F0781F80FFC000000007FE03F07C3C3871C639CCE66666CD936DB6DA5A";
defparam ram_block1a52.mem_init1 = "5AD4AD56AAA55552AAB55A95A52D25B6DB24C99B33399CE738E3C78787C0FE007FFFFFFFFE00FE07C3E3C38E39CE733999B326C9B6DB4B4B4A56AD54AAAAAAAAB55AB5294B4B6924DB264CCCCCCE739C71C78787C0FC03FFF8000FFFE01FC1F0F0F1C71C633999C999B26D924B69694A56A9552AAAAAA555AB52B4A5B49249364CD9999CCE738E3870F0F83F807FFE0000FFFC03F03E1E1C38E31CC66333266CDB2492DA5AD6B56AB5555555554AA54A5296D25B649B36666666339C71C78F0F83F01FF800000007FE03F07C3C38F38E7399CCCD99324DB6D25A5294A954AAAAAAAAA954AD4A5ADA49249366CCCCCCE631C71C78F87C1FC01FFFFFFFFFC01FC1";
defparam ram_block1a52.mem_init0 = "F0F8F1C71C633999999326C92492D2D6B52A556AAAAAAA955AB5294B496DB6499336667339CE39E38787C1F807FFC00001FFF01F81E0F1E38E31CC6666666CDB24925A5A5295AAD554AAAD555AA56A52D2DB6DB64D99333399CE31C70E1E0F81FC007FFFFFFC007F03E0F0E1C718E63399993364DB6DB496B5AD5AA5555555555AAD4AD69692DB649B3666666339C638F1E1E0FC07F8000000000FF81F83C3C78E39CE73333332649B6DB4B4B5AD5AA55556A55552A95A96B496DB6D93666CCE66318E38E1C3E1F81FF00007F00007F80F83C3C38E39CE733333326C9B6DA4B4A52952AB555555552AB56B5AD2DA4936C9933333318C638E3C3C3E0FE01FFFFF";

cyclonev_ram_block ram_block1a76(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a76_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a76.clk0_core_clock_enable = "ena0";
defparam ram_block1a76.clk0_input_clock_enable = "ena0";
defparam ram_block1a76.clk0_output_clock_enable = "ena0";
defparam ram_block1a76.data_interleave_offset_in_bits = 1;
defparam ram_block1a76.data_interleave_width_in_bits = 1;
defparam ram_block1a76.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a76.init_file_layout = "port_a";
defparam ram_block1a76.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a76.operation_mode = "rom";
defparam ram_block1a76.port_a_address_clear = "none";
defparam ram_block1a76.port_a_address_width = 13;
defparam ram_block1a76.port_a_data_out_clear = "none";
defparam ram_block1a76.port_a_data_out_clock = "clock0";
defparam ram_block1a76.port_a_data_width = 1;
defparam ram_block1a76.port_a_first_address = 24576;
defparam ram_block1a76.port_a_first_bit_number = 4;
defparam ram_block1a76.port_a_last_address = 32767;
defparam ram_block1a76.port_a_logical_ram_depth = 65536;
defparam ram_block1a76.port_a_logical_ram_width = 24;
defparam ram_block1a76.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a76.ram_block_type = "auto";
defparam ram_block1a76.mem_init3 = "1E1C3C3C7878F0F1E1E1C3C3C787870F0F0E1E1E1C3C3C3C3C78787878787878787878787878787C3C3C3E1E1E0F0F8783C3E1E0F0783C1E0F07C3E0F07C1F0F83E0F83E0F81F07C0F83F07E0FC0F81F81F81F81F80FC07E03F01FC07F80FF01FE01FE00FF007FC00FF800FFC007FF8007FFE0007FFF80000FFFFF80000003FFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFF80003FFF8003FFC007FF007FE00FF00FF00FE03F80FC07E07E07C0F81F07C1F07C3E1F0F8783C3C3C3C3C7870F1E3C78E1C78E3871C71C71C638E31C639C631CE739CE7319CE673198CCE66733331999999999933332666CC99B3264D9B26C9B26C936C936DB6492492496DB69";
defparam ram_block1a76.mem_init2 = "25B496D2D25A5A5A52D294B5AD6B5A94AD4AD5AB56AD52A954AAD552AA95555AAAAAAAA5555556AAAAAAA95554AAA555AA954AB54A952B52B52B5AD6B5A52D696969692D25B6925B6DB6DB6D924DB26D9366C993266CCC99999933999999CCC663398CE739CE31CE38C71C71E38F1C3C7870F0F8783C1F07C0FC0FC07F00FF003FF8003FFFFE000000000001FFFFE0007FF007FC07F01F81F03E0F87C3C3C3C3C78F1C38E38E39C738C6318C673199CCCC666666CCCD99B366C9B26C926DB6DB6DB692DA4B4B4B4A5AD6B5295AB56AD56AB554AAAB555555555555552AAAD55AA956AD5A95A94A5296B4B4B496D24B6DB6DB249B26C9B366CCD9999999998CCE";
defparam ram_block1a76.mem_init1 = "6339CE738C71CE3871C3870F0F0F0783E0FC0FC03F803FF8000FFFFFFFFFFFFFE0003FF007F80FC0FC1F0783C3C3C78F1C71C71C639CE7319CCE6666666664CC99364D936DB2492DB496D2D2D296B5295A956A954AAB55556AAAAAAB55556AA954AB56A56A5296B4B4B496DA49249B6C9B26CD9B3332663333198CE739C638E38E3870E1E1F0F83E0FC07F807FF0001FFFFFFFFFE0003FF807F81F81F0783C3C3870E38E38E718C673199CCCCCCD99B366C9B64924924B692D2D294A52B52A55AA95552AAAAAAAAA9555AA956AD5A94A52D2D2D25B6DB6DB24D93264CCC999CCCC67318C738E38E3870F0F0F83E0FC07F803FFE000000000003FFC00FE03F07E";
defparam ram_block1a76.mem_init0 = "1F0F0F1E3C71C738C7318CC666666664CD9324DB24924B692D2D694A56AD5AA554AAAAAAAAAAAAAD55AA55A95AD694B496924B64926C9B3664CCCCCCE67318C738E38E3C78787C3E07E03FC00FFFFC00001FFFF801FE03F07E1F0F0E1C38E38C739CC66733333266CD9364924924B69694B5A95A956AA55552AAAAB5555AA956AD4A52D69692DB6DB6C9366CD99999998CC6318E71C70E1C3C3E0F81F807FE0003FFFFFF0001FF807E07C1E0F1E1C71C71CE7399CCCCCCCC99326D924925B49694A5295AA55AAAD55555555AAAD56AD4AD694B496D24924D9364CC999998CC6738C71C71E3C3C3E0FC0FE00FFFC0000001FFF803F81F83E1E1E3C71C738C6731";

cyclonev_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 8191;
defparam ram_block1a4.port_a_logical_ram_depth = 65536;
defparam ram_block1a4.port_a_logical_ram_width = 24;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init3 = "19CC639C71C78F0F0F83F03F803FFF00000007FFE00FE07E0F87878F1C71C639CC66333332664D936492496D25A52D6A56AD56AAB555555556AAB54AB5294A52D25B4924936C993266666667339CE71C71C70F1E0F07C0FC03FF0001FFFFFF8000FFC03F03E0F87870E1C71CE318C663333333366CD926DB6DB692D2D694A56AD52AB5555AAAAA95554AAD52B52B5A52D2DA4924924D9366CC999999CCC6739C638E3870E1E1F0FC1F80FF003FFFF000007FFFE007F80FC0F87C3C3C78E38E39C6319CCE6666664CD9B26C924DA492D25A52D6B52B54AB556AAAAAAAAAAAAA554AB56AD4A52D69692DA49249B64993664CCCCCCCC66319C639C71C78F1E1E1F0";
defparam ram_block1a4.mem_init2 = "FC1F80FE007FF800000000000FFF803FC07E0F83E1E1E1C38E38E39C6319CC66673326664C993649B6DB6DB496969694A52B56AD52AB5552AAAAAAAAA95552AB54A95A94A52969692DA4924924DB26CD9B3366666673319CC631CE38E38E1C3878783C1F03F03FC03FF8000FFFFFFFFFF0001FFC03FC07E0F83E1F0F0E1C38E38E38C739CE63319998CC9999B366C9B26DB24924B6D25A5A5AD294AD4AD5AA552AAD5555AAAAAAAD5555AAA552AD52B5295AD2969696D25B69249B6D9364D932664CCCCCCCCCE67319CE738C71C71C71E3C7878783C1F07E07E03FC01FF8000FFFFFFFFFFFFFE0003FF803F807E07E0F83C1E1E1E1C3871C38E71C639CE7398C";
defparam ram_block1a4.mem_init1 = "E663333333333666CD9B26C9B249B6DB6DA496D25A5A5AD294A52B52B56AD52AB556AAA955555555555555AAAA555AAD56AD5AB5295AD6B4A5A5A5A4B692DB6DB6DB6C926C9B26CD9B336666CCCCCC66673319CC6318C639C738E38E3871E3C787878787C3E0F81F03F01FC07FC01FFC000FFFFF000000000000FFFFF8003FF801FE01FC07E07E07C1F0783C3E1E1C3C7871E38F1C71C638E718E739CE63398CC66733333399333332666CC99326CD936C9B64936DB6DB6DB492DB49692D2D2D2D694B5AD6B5A95A95A952A55AA552AB554AAA55552AAAAAAAD555554AAAAAAAB55552AA9556AA552A956AD5AB56A56A52B5AD6B5A529694B4B4B49696D25B49";
defparam ram_block1a4.mem_init0 = "2DB6D24924924DB6D926D926C9B26C9B364C99B3266CCC99999333333333319999CCCE663319CCE7319CE739CE718C738C718E38C71C71C71C38E3C70E3C78F1E1C3C78787878783C3E1F0F87C1F07C1F03E07C0FC0FC07E03F80FE01FE01FE00FFC01FFC007FF8003FFF80003FFFFE0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFF80000003FFFFE00003FFFC000FFFC003FFC007FE003FE007FC01FE00FF00FF01FE03FC07F01F80FC07E03F03F03F03F03E07E0FC1F83E07C1F03E0F83E0F83E1F07C1E0F87C1E0F0783C1E0F0F8783C3E1E0F0F0F878787C3C3C3C3C3C3C3C3C3C3C3C3C3C3C7878787870F0F0E1E1E1C3C3C787870F0F1E1E3C3C787870F0";

cyclonev_ram_block ram_block1a28(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.clk0_output_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "rom";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "clock0";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 8192;
defparam ram_block1a28.port_a_first_bit_number = 4;
defparam ram_block1a28.port_a_last_address = 16383;
defparam ram_block1a28.port_a_logical_ram_depth = 65536;
defparam ram_block1a28.port_a_logical_ram_width = 24;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init3 = "FFFFF00FE0F87878E38C631999999326D924B696B5AD5AA955555555AA95294A5A4B6DB26C9999999CE738E3878783E03FC0001FC0001FF03F0F870E38E318CCE66CCD936DB6D25AD2B52A95554AD5554AB56B5A5A5B6DB24C9999999CE738E3C78783F03FE0000000003FC07E0F0F1E38C7398CCCCCD9B24DB692D2D6A56AB5555555554AB56B5AD25B6DB64D99333398CE31C70E1E0F81FC007FFFFFFC007F03E0F0E1C718E73399993364DB6DB69694AD4AB5556AAA5556AB5294B4B49249B66CCCCCCC6718E38F1E0F03F01FFF000007FFC03F07C3C38F38E7399CCCD99324DB6D25A5295AB552AAAAAAAD54A95AD696924926C9933333398C71C71E3E1F";
defparam ram_block1a28.mem_init2 = "07F007FFFFFFFFF007F07C3E3C71C718CE666666CD924924B6B4A56A552AAAAAAAAA552A5294B496DB6499336667339CE39E38787C1F80FFC00000003FF01F83E1E3C71C7398CCCCCCD9B24DB496D294A54AA5555555555AAD5AD6B4B69249B66CC9998CC6718E3870F0F81F807FFE0000FFFC03F83E1E1C38E39CE673333664D924925B4A5A95AB554AAAAAA9552AD4A52D2DA4936C9B332733398C71C71E1E1F07F00FFFE0003FFF807E07C3C3C71C739CE6666664C9B6492DA5A5295AB55AAAAAAAAA556AD4A5A5A5B6DB26C99B33399CE738E3878F87C0FE00FFFFFFFFFC00FE07C3C3C78E39CE733999B32649B6DB49694B52B55AAA95554AAAD56A56B4";
defparam ram_block1a28.mem_init1 = "B4B6DB6D9366CCCCCE6738C71C38787C1F80FFC000000007FE03F03C1E3C71C718C667333664C936DB692D296A56A9556AAAAAA555AA56A52D2DA49249B266CCCCC66318E38E1C3C3E07E01FFC0000001FFE03F83E1E1E38638C631999999B364DB6DB49694B52B54AAB5555556AA956A56B4B4B6924DB26CC99998CC6318E38F1E1F0FC0FE003FFFFFFFF801FE07C1F0E1C38E718C663333366CDB24924B4B4B52952A95552AAAD555AAD5A94B5A4B6DB6D9366CCCCCCC6738C71C78F0F87E07F003FFFFFFFFFC00FE07C1E0E1C38E31CC6733333366CDB2492DA4B5A56A54AA55555555555AAD5295A52D25B6DB64D93326663339CE71C71E3C3C1F03F807F";
defparam ram_block1a28.mem_init0 = "FF00000FFFE01FC0F83C3C78E38E719CC666666CD9B6492496D2D294AD5AA5556AAAAA9555AA54AD694B496DB6D9264C9999998CE639C71C78F0F07C0FC01FFE00000003FFC03F83E0F0F0E1C718E7399CCCCCC99324DB6DB692D296A56AD52AAB555555AAAD56AD4A52D2D2DB6DB64D9336666673398E71C71C38787C1F81FE007FFFFFFFFFC00FF01F07C3C3C78E39C6318CCC666CCD9B24DB6DB4969694AD4A956AAB5555555AAAD56AD4A52D6D2DB4936D9366CCCCCCCC6739CE38E3878F0783F03FC01FFFF0000FFFF803FC0FC1E0F0E1C71C718C673399999B326C9B6492DB4B4B4A56B56AB556AAAAAAAAAD55AA54AD6B5A5A4B6D26DB26C993333333";

cyclonev_ram_block ram_block1a101(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a101_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a101.clk0_core_clock_enable = "ena0";
defparam ram_block1a101.clk0_input_clock_enable = "ena0";
defparam ram_block1a101.clk0_output_clock_enable = "ena0";
defparam ram_block1a101.data_interleave_offset_in_bits = 1;
defparam ram_block1a101.data_interleave_width_in_bits = 1;
defparam ram_block1a101.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a101.init_file_layout = "port_a";
defparam ram_block1a101.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a101.operation_mode = "rom";
defparam ram_block1a101.port_a_address_clear = "none";
defparam ram_block1a101.port_a_address_width = 13;
defparam ram_block1a101.port_a_data_out_clear = "none";
defparam ram_block1a101.port_a_data_out_clock = "clock0";
defparam ram_block1a101.port_a_data_width = 1;
defparam ram_block1a101.port_a_first_address = 32768;
defparam ram_block1a101.port_a_first_bit_number = 5;
defparam ram_block1a101.port_a_last_address = 40959;
defparam ram_block1a101.port_a_logical_ram_depth = 65536;
defparam ram_block1a101.port_a_logical_ram_width = 24;
defparam ram_block1a101.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a101.ram_block_type = "auto";
defparam ram_block1a101.mem_init3 = "783E0F83F03F80FF007FF0003FFFFF8000000FFFFFE0007FF007F80FE07E07C1F0F87C3C3878F1E38F1C718E39CE318C673198CCC66666666CCCD99326CD936C936D92492DB6925A4B4B4B4A5AD6B5A95A952A55AA554AAB5555AAAAAAAAAAAAAA55552AA955AAD5AA56AD4A56B5A52D6969696D25B6924924924DB64DB264D9B3666CCCCD9999CCCCE663398CE739C631C738E38E1C70E1C3C78787C3E1F07C0F81FC0FF01FF003FF8000FFFFFFFC0001FFFFFFF0000FFE007FC03F80FC0FC1F83E1F0F8787870F1E3C71E38E38E71CE31CE7398C6733998CCCCCCCCCCCCD99B3264C9B26C9B249B6D92496DB6925B4B6969696B4A5AD6B5295A952A54AB55A";
defparam ram_block1a101.mem_init2 = "A9552AAA555556AAAAAAAAAAB555556AAA555AA954AB56AD5A95A94AD6B4A5AD2D2D2D2DA5B6925B6DB6DB6D924DB26D9326CD9B3666CCCD999999999CCCC667319CC6739CE318E71C638E38E3C71E3C78F0E1E1E1F0F87C1F07C1F81F81FC07F807FC007FF0003FFFFC00000000000000003FFFFC000FFF003FE00FE01F80FC0FC0F83E0F83C1E1E1E1E1E1C3870E3C71C78E39C71CE39C6318C6318CE633998CCE6666733333266666CCC99B366CD9326C9B64DB249B6DB6CB6DB6DA496D25B4B696969696B4A5AD6B5AD4A56A56A54A952AD52A955AAB554AAA955556AAAAAAAAAAAAAAAAAAAAD55552AAA5552AA556AB54AB54A952B52B52B5294A5294A5";
defparam ram_block1a101.mem_init1 = "AD2D696969696D2DA4B6925B6D24924924924DB64936C9B64D9366C993264CD993326666CCCCCCCCCCCCCC666733399CCE63398C6739CE738C639C738E71C71C71C71C70E3871E3C78F0E1E1E3C3C1E1E0F0783C1F07C1F83F07E07E03F01FC07F807F803FE003FF8007FFC0003FFFFE000000003FFFFFFFFFFC000000003FFFFC0001FFF8007FF001FF003FC03FC03F80FE03F03F81F03F07E0F83E0F83C1F0F8783C3C3C3C3C3C3C7870E1E3870E3C70E38F1C71C71C71C71CE38C718E31CE318E739CE739CE6319CC67319CCE6733998CCCE6667333333333999B3333333326666CCC999B32664C99B366CD9B364D9B26C9B26C9B64DB26D924DB24936DB2";
defparam ram_block1a101.mem_init0 = "4924936DB6DB4924924B6DA492DB492DA4B692DA4B49696D2D2DA5A5A5A5AD2D2D696B4A5AD296B5A5294A5294A52B5AD4A56B52B5A95A95AB52B56A54A952A54A956A952AD52A956AB55AAD56AA556AAD55AAB556AAB555AAAD555AAAB5555AAAA955554AAAAA95555556AAAAAAAAA555555555555555555555555555555555555555555AAAAAAAAAAD5555554AAAAAAD55555AAAAAD5555AAAA95554AAAA5554AAA9555AAA9555AAAD552AA9556AA9552AAD55AAB556AA554AAD54AA955AAD54AAD56AA552A954AA556A954AA552A956AB54AA55AAD52AD52A956A956A956A956A956A956AD52AD52AD5AA55AB54AB56A956AD52A55AB54AB56A952AD5AA54";

cyclonev_ram_block ram_block1a125(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a125_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a125.clk0_core_clock_enable = "ena0";
defparam ram_block1a125.clk0_input_clock_enable = "ena0";
defparam ram_block1a125.clk0_output_clock_enable = "ena0";
defparam ram_block1a125.data_interleave_offset_in_bits = 1;
defparam ram_block1a125.data_interleave_width_in_bits = 1;
defparam ram_block1a125.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a125.init_file_layout = "port_a";
defparam ram_block1a125.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a125.operation_mode = "rom";
defparam ram_block1a125.port_a_address_clear = "none";
defparam ram_block1a125.port_a_address_width = 13;
defparam ram_block1a125.port_a_data_out_clear = "none";
defparam ram_block1a125.port_a_data_out_clock = "clock0";
defparam ram_block1a125.port_a_data_width = 1;
defparam ram_block1a125.port_a_first_address = 40960;
defparam ram_block1a125.port_a_first_bit_number = 5;
defparam ram_block1a125.port_a_last_address = 49151;
defparam ram_block1a125.port_a_logical_ram_depth = 65536;
defparam ram_block1a125.port_a_logical_ram_width = 24;
defparam ram_block1a125.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a125.ram_block_type = "auto";
defparam ram_block1a125.mem_init3 = "0000000FFF007F80FC1F83C1E1E1E3C71C39C718C6319CCE66666666CC99326C926DB6DB496D2D2D294A52B56AD52AB5554AAAAAAAAAB5556AA55AA56A52B4A5A5A5A4B6DB6DB649B26CD9B333333333198CE739C638E38E1C3878787C1F07E03F803FF0000FFFFFFFFF80007FE00FE03E07C1F0F0F0E1C38E38E31CE7398CC6666666664CD9B26C936DB6DB692D25A52D6B5A952A55AAD554AAAAAAAAAAAA5556AB54A952B5AD694B4B692DB6DB6DB26C9B266CCCC998CCCE67318C738E71C78E1C3C3C3C1F07E07F00FF800FFFFF80000FFFFF8007FC07F03F07C1E0F0E1E3871C71CE31CE633998CCCCCCC999326C9B249B6DB492DA5A5A5294A56A54AB55";
defparam ram_block1a125.mem_init2 = "AAAD5555555555555AAAD56A952B5294A52D2D2DA496DB6D926D93264CD999999999CCE7318C718E38E3C70F1E0F0F83E07E07F803FF80001FFFFFFF80001FFC01FC07E07C1F0F0F0F1E3C71C718E718CE73399999999993366C9B26DB6496DB49692D696B5AD4AD5AA552AAD555552AA9555556AA954AB56A56B5AD29696D25B6924936C9364C9933366666633319CC631CE38C70E3870F0F0F07C1F03F01FE00FFF0000007FE000000FFF803FC07E07C1F078787870E38F18E39C6319CC66333333332664C9B26C936DB6DB492D2DAD2D6B5AD4A952AD54AAA55555555555554AAA556A952A56B5AD696B696925B6DB6DB24D9366CC99993331999CCE6318C";
defparam ram_block1a125.mem_init1 = "738E38E38F1E3C3C3E1F07E0FE07F803FF80001FFFFFFFF00003FF803FC07E07C0F0783C3878E1C71C71CE318C6733998CCCCCD9993264D9364936DB6925B49696B4A5A94AD4A956AB554AAAAB5555556AAAA9556AB54A95A95AD694B4B4B692DB6DB6DB24D9366CC999B33333199CCE6318C738E31E38E1C3C787C3C1F03E07F01FF003FFF00000000000001FFF801FE01F80F81F0787C3C3870E3C71C638C739CC63319998CCD99993366C9B26D924924925B4969696B4A5295A952AD52AB5552AAAAAAAAAAAAAB5552AB54AB52A52B5AD2969696D25B6D249B6C9364D932664CCCCCCCCCC663398C631C638E38E3C78F0E1F0F07C1F03F01FC01FF8007FFF";
defparam ram_block1a125.mem_init0 = "FFC0003FFFFFE001FF803F80FC0F83E0F0787870E1C78E38E71CE719CE6331998CCCCC99993364C9B26DB24924925B692D2D2D294A5295A952A552A9554AAAAA55555552AAAA9556AA55AA56AD6A5294B5A5A5B4B6D24924924DB24D93264CD999333331999CCE6339CE31CE38E38E3C78F1E1E1F0F83E0FC0FC07F803FF8001FFFFFFFFFFFFFFF0003FF803FC07F03E07C1E0F0F8F0F1E3871C71C718E739CE73198CCCE666666CCC99B364C9B649B6DB6DB6DA4B696969694A5294AD4A952AD56AA5556AAAAAAB552AAAAAA9555AA954AB56AD4AD6A52D694B4B496D25B6DB6DB6D926C9B26CD9933266666666633399CC6318C639C71C71C71E3878F0F0F0";

cyclonev_ram_block ram_block1a149(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a149_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a149.clk0_core_clock_enable = "ena0";
defparam ram_block1a149.clk0_input_clock_enable = "ena0";
defparam ram_block1a149.clk0_output_clock_enable = "ena0";
defparam ram_block1a149.data_interleave_offset_in_bits = 1;
defparam ram_block1a149.data_interleave_width_in_bits = 1;
defparam ram_block1a149.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a149.init_file_layout = "port_a";
defparam ram_block1a149.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a149.operation_mode = "rom";
defparam ram_block1a149.port_a_address_clear = "none";
defparam ram_block1a149.port_a_address_width = 13;
defparam ram_block1a149.port_a_data_out_clear = "none";
defparam ram_block1a149.port_a_data_out_clock = "clock0";
defparam ram_block1a149.port_a_data_width = 1;
defparam ram_block1a149.port_a_first_address = 49152;
defparam ram_block1a149.port_a_first_bit_number = 5;
defparam ram_block1a149.port_a_last_address = 57343;
defparam ram_block1a149.port_a_logical_ram_depth = 65536;
defparam ram_block1a149.port_a_logical_ram_width = 24;
defparam ram_block1a149.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a149.ram_block_type = "auto";
defparam ram_block1a149.mem_init3 = "1E1E1E3C38F1C71C71C738C6318C6733998CCCCCCCCC9993366C9B26C936DB6DB6DB496D25A5A52D694AD6A56AD5AA552AB5552AAAAAA955AAAAAAAD554AAD56A952A56A5294A52D2D2D2DA4B6DB6DB6DB24DB264D9B32666CCCCCCE6663319CE739CE31C71C71C38F1E1E3E1E0F07C0F81FC07F803FF8001FFFFFFFFFFFFFFF0003FF803FC07E07E0F83E1F0F0F1E3C78E38E38E718E7398CE67333199999333664C993649B6492492496DA5B4B4B5A5294AD6AD4AB54AAD552AAAA95555554AAAAA5552A954A952B5294A5296969692DB49249249B6C9B264D99333266666333198CE731CE71CE38E3C70E1C3C3C1E0F83E07E03F803FF000FFFFFF80007FF";
defparam ram_block1a149.mem_init2 = "FFFC003FF007F01F81F07C1E1F0E1E3C78E38E38C718C63398CC66666666664CC99364D926DB2496DB496D2D2D296B5A94A95AA55AA9555AAAAAAAAAAAAAA9555AA956A952B5294A5AD2D2D25B4924924936C9B26CD9933336663333198C6739C638C71C78E1C38787C3C1F03E03F00FF003FFF00000000000001FFF801FF01FC0F81F0787C3C7870E38F18E39C6318CE6733199999B33266CD93649B6DB6DB692DA5A5A52D6B52B52A55AAD552AAAAD555555AAAAA555AAD52A56A52B4A5AD2D25B492DB6D924D9364C9933366666633399CC6318E71C71C70E3C38783C1E07C0FC07F803FF80001FFFFFFFF00003FF803FC0FE0FC1F0F87878F1E38E38E39C";
defparam ram_block1a149.mem_init1 = "6318CE673331999333266CD93649B6DB6DB492D2DAD2D6B5AD4A952AD54AAA55555555555554AAA556A952A56B5AD696B696925B6DB6D926C9B264CC999999998CC67318C738E31E38E1C3C3C3C1F07C0FC07F803FFE000000FFC000001FFE00FF01F81F07C1E1E1E1C38E1C638E718C6731998CCCCCD9993264D926D92492DB496D2D296B5AD4AD5AA552AAD555552AA9555556AA954AB56A56B5AD2D692D25B6D24DB6C9B26CD99333333333399CE631CE31C71C78F1E1E1E1F07C0FC07F007FF00003FFFFFFF00003FF803FC0FC0F83E1E0F1E1C78E38E31C6319CE67333333333664C9936C936DB6D24B6969694A5295A952AD56AAB55555555555556AAB";
defparam ram_block1a149.mem_init0 = "55AA54AD4A5294B4B4B6925B6DB249B26C99332666666633398CE718E71C71C38F0E1E0F07C1F81FC07FC003FFFFE00003FFFFE003FE01FC0FC1F078787870E3C71CE39C6319CCE6663326666CC9B26C9B6DB6DB692DA5A52D6B5A952A55AAD554AAAAAAAAAAAA5556AB54A952B5AD694B49692DB6DB6D926C9B3664CCCCCCCCC66339CE718E38E3870E1E1E1F07C0F80FE00FFC0003FFFFFFFFE0001FF803F80FC1F07C3C3C3870E38E38C739CE6331999999999B366C9B24DB6DB6DA4B4B4B4A5A94AD4AB54AAD555AAAAAAAAAA5555AA956AD5A94A52969696D25B6DB6C926C993266CCCCCCCCE67318C631C73871C78F0F0F0783F07E03FC01FFE0000000";

cyclonev_ram_block ram_block1a173(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a173_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a173.clk0_core_clock_enable = "ena0";
defparam ram_block1a173.clk0_input_clock_enable = "ena0";
defparam ram_block1a173.clk0_output_clock_enable = "ena0";
defparam ram_block1a173.data_interleave_offset_in_bits = 1;
defparam ram_block1a173.data_interleave_width_in_bits = 1;
defparam ram_block1a173.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a173.init_file_layout = "port_a";
defparam ram_block1a173.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a173.operation_mode = "rom";
defparam ram_block1a173.port_a_address_clear = "none";
defparam ram_block1a173.port_a_address_width = 13;
defparam ram_block1a173.port_a_data_out_clear = "none";
defparam ram_block1a173.port_a_data_out_clock = "clock0";
defparam ram_block1a173.port_a_data_width = 1;
defparam ram_block1a173.port_a_first_address = 57344;
defparam ram_block1a173.port_a_first_bit_number = 5;
defparam ram_block1a173.port_a_last_address = 65535;
defparam ram_block1a173.port_a_logical_ram_depth = 65536;
defparam ram_block1a173.port_a_logical_ram_width = 24;
defparam ram_block1a173.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a173.ram_block_type = "auto";
defparam ram_block1a173.mem_init3 = "54AB56A952AD5AA55AB54A956AD52AD5AA55AB54AB56A956A956AD52AD52AD52AD52AD52AD52A956A956AB54AA55AAD52A954AA552AD54AA552A954AAD56AA556AB552AA556AA554AAD55AAB556AA9552AAD552AA9556AAB5552AAB5552AAA5554AAAA55552AAAB55556AAAAB555556AAAAAA55555556AAAAAAAAAB555555555555555555555555555555555555555554AAAAAAAAAD5555552AAAAA555552AAAB5555AAAB5556AAB555AAAD55AAB556AAD54AAD56AB55AAD52A956A952AD52A54A952A54AD5A95AB52B52B5A95AD4A56B5A94A5294A5294B5AD296B4A5AD2D69696B4B4B4B4B69696D2D25A4B692DA4B6925B6924B6DA4924925B6DB6D924924";
defparam ram_block1a173.mem_init2 = "9B6D9249B64936C9B64DB26C9B26C9B364D9B366CD9B3264CC99B332666CCCC999999999B333999999999CCCCE66633399CCE67319CC67318CE739CE739CE318E718E31C638E71C71C71C71C71E38E1C78E1C38F0E1C3C787878787878783C3E1F0783E0F83E0FC1F81F03F81F80FE03F807F807F801FF001FFC003FFF00007FFFF8000000007FFFFFFFFFF800000000FFFFF80007FFC003FF800FF803FC03FC07F01F80FC0FC1F83F07C1F0783C1E0F0F07878F0F0E1E3C78F1C38E1C71C71C71C71CE39C738C639CE739CC63398CE6733999CCCC66666666666666CCCC99933664C99326CD9364DB26D924DB6492492492496DB492DA4B696D2D2D2D2D696B";
defparam ram_block1a173.mem_init1 = "4A5294A5295A95A95A952A55AA55AAD54AA9554AAA955556AAAAAAAAAAAAAAAAAAAAD55552AAA555AAB552A956A952A54AD4AD4A56B5AD6B4A5AD2D2D2D2DA5B496D24B6DB6DA6DB6DB249B64DB26C99366CD9B32666CCCCC999999CCCCCE6633398CE6318C6318C738E71C738E3C71C78E1C3870F0F0F0F0F0783E0F83E07E07E03F00FE00FF801FFE0007FFFF800000000000000007FFFF8001FFC007FC03FC07F03F03F07C1F07C3E1F0F0F0E1E3C78F1C78E38E38C71CE318E739CC67319CCC66673333333336666CCD9B366C9936C9B64936DB6DB6DB492DB4B696969696B4A5AD6A52B52B56AD5AA552AB554AAAD55555AAAAAAAAAAAD55554AAA9552A";
defparam ram_block1a173.mem_init0 = "B55AA54A952B5295AD6B4A5AD2D2D2DA5B492DB6D24936DB249B26C9B264C99B33666666666666633399CC6339CE718E71CE38E38F1C78F1E1C3C3C3E1F0F83F07E07E03F807FC00FFE0001FFFFFFF00007FFFFFFE0003FF801FF01FE07F03E07C1F0F87C3C3C7870E1C70E38E39C718C739CE63398CCE6667333366666CCD9B364C9B64DB6492492492DB496D2D2D2D694B5AD4A56AD4AB56AB552AA95554AAAAAAAAAAAAAB5555AAA554AB54A952B52B5AD6B4A5A5A5A4B492DB6924936D926D9366C99336666CCCCCCCC6663319CC6318E738E31C71E38F1E3C38787C3E1F07C0FC0FE03FC01FFC000FFFFFE0000003FFFFF8001FFC01FE03F81F83E0F83C";

cyclonev_ram_block ram_block1a53(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a53_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a53.clk0_core_clock_enable = "ena0";
defparam ram_block1a53.clk0_input_clock_enable = "ena0";
defparam ram_block1a53.clk0_output_clock_enable = "ena0";
defparam ram_block1a53.data_interleave_offset_in_bits = 1;
defparam ram_block1a53.data_interleave_width_in_bits = 1;
defparam ram_block1a53.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a53.init_file_layout = "port_a";
defparam ram_block1a53.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a53.operation_mode = "rom";
defparam ram_block1a53.port_a_address_clear = "none";
defparam ram_block1a53.port_a_address_width = 13;
defparam ram_block1a53.port_a_data_out_clear = "none";
defparam ram_block1a53.port_a_data_out_clock = "clock0";
defparam ram_block1a53.port_a_data_width = 1;
defparam ram_block1a53.port_a_first_address = 16384;
defparam ram_block1a53.port_a_first_bit_number = 5;
defparam ram_block1a53.port_a_last_address = 24575;
defparam ram_block1a53.port_a_logical_ram_depth = 65536;
defparam ram_block1a53.port_a_logical_ram_width = 24;
defparam ram_block1a53.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a53.ram_block_type = "auto";
defparam ram_block1a53.mem_init3 = "E1E1E1E3C70E38F18E38C739CE7398CC667333333333666CC99366C936C924DB6924B6D2DA5A5AD296B5A95A95AB54AA554AAAD555554AAAB5555552AAB556AB56A95A95AD6B5AD2D2D2D25B4924B6C924DB24D93264CD9993333333999CCE6319CE31CE38E38E3870E1E3C3E1E0F83F07E03F807FC00FFFE000000000000000FFFC007FC03F81F81F03C1E0F0F0E1E3871C71C718E718C673198CCC666666CCCD9B366C9B24DB6DB6DB6D25B4B4B4A5AD6B5A95AB54AB552AAD55552AAAAAAA555552AAD54AB56AD4AD6A5AD6969696D25B6DB6DB6C9364D93266CCC999999CCCC67319CE718E31C71C38F1E3C3C3C1F0FC1F81FC07F801FFF000001FFFFE00";
defparam ram_block1a53.mem_init2 = "0003FFE007F80FE07E0F83E1F0F0E1E3871C71C718E739CE6733999999999993366C9926C924DB6D24B692D2D2D694A52B52A54AA556AAB555555555555554AAA556AB56AD4AD6B5AD2D2D2DA4B6DB6DB6D936C993266CCCD9998CCCE67318C639C638E3871E3C78787C3E0FC1F80FE00FFC000FFFFFFFFFFFFFF0007FE00FE03F03E0F87C3C3C78F1C78E31C639CE7319CCCE666666CCC99326C9B6492492496D25A5A5A5294AD6AD5AA552AAD5555AAAAAAAD5555AAA552AD5A95A94A5AD2D2DA5B6924926DB24D9B266CCD999999CCCE6339CE718E38E38E1C3C787C3C1F03F03F80FF8007FFFC000000007FFFC007FC03F81F83E0F0787870E1C71C71C63";
defparam ram_block1a53.mem_init1 = "9CE73198CCC66664CCD99326C9B6492492496D2DA5AD294A52B56AD52A9554AAAAAAAAAAAAAA5552A956A95A94A5296B4B696DA4924926D926CD9B326666666673398CE738C718E3C71E3C3C3C3E0F83F03F807FC003FFFFF8000FFFFFE001FF00FE07E07C3E1E0E1E3C71E38C718E7398CE663333333666CD9B26C926DB6DA49692D2D694A52B52A55AAD552AAAAB5555AAAAA9556AB54A95A94A52D69692DA496DB649364D93266CCCCCCCCCC66339CE71CE38E3870E1E1E1E0F83F03F80FF800FFFF800000007FFFC007FC03F03F07C1E0F0E1E3C71C71C639CE73198CCCCCCCCCD99366C936C924925B4969696B4A56A56AD52A9556AAAAAAAAAAAAAB554";
defparam ram_block1a53.mem_init0 = "AA55AB52B5296B4B4B496DA49249B64D9366CCD99999998CC67318C738E38E3870F1E1F0F83E07E07F803FF800003FFFFE00001FFE00FE03F03E0F8787878F1C38E39C639CE6331998CCC99993364C9B6492492496D25A5AD294A56A54AB552AA95555555555552AA955AA54AD4A5296B4B496D24924924D9364C99333333333399CC6318E71C71C78F1E1E1E0F83E07F01FE003FFF8000000000FFFE003FC07F03E0F83C3C3C3871C71C738C6319CC66667366664CD9324D924924925B4B694B4A52B52B56AB552AAA55555555552AAA556A956A56B5AD6969696DA4924926D9364C99933333333198CE739CE39C70E3870F0F0F07C1F81FC03FE001FFFFFFF";

cyclonev_ram_block ram_block1a77(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a77_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a77.clk0_core_clock_enable = "ena0";
defparam ram_block1a77.clk0_input_clock_enable = "ena0";
defparam ram_block1a77.clk0_output_clock_enable = "ena0";
defparam ram_block1a77.data_interleave_offset_in_bits = 1;
defparam ram_block1a77.data_interleave_width_in_bits = 1;
defparam ram_block1a77.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a77.init_file_layout = "port_a";
defparam ram_block1a77.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a77.operation_mode = "rom";
defparam ram_block1a77.port_a_address_clear = "none";
defparam ram_block1a77.port_a_address_width = 13;
defparam ram_block1a77.port_a_data_out_clear = "none";
defparam ram_block1a77.port_a_data_out_clock = "clock0";
defparam ram_block1a77.port_a_data_width = 1;
defparam ram_block1a77.port_a_first_address = 24576;
defparam ram_block1a77.port_a_first_bit_number = 5;
defparam ram_block1a77.port_a_last_address = 32767;
defparam ram_block1a77.port_a_logical_ram_depth = 65536;
defparam ram_block1a77.port_a_logical_ram_width = 24;
defparam ram_block1a77.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a77.ram_block_type = "auto";
defparam ram_block1a77.mem_init3 = "AB56A956AD52A55AB54A956A952AD5AA55AB54AB56A956A956AD52AD52AD52AD52AD52AD52AD52A956A954AB54AA552AD56AB54AA552A954AA556AB55AA955AAD54AAD54AAD55AA9552AA554AA9552AAD552AAD552AA9554AAA5556AAAD555AAAB5554AAAA55556AAAAD55556AAAAAD555554AAAAAAAD5555555552AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5555555556AAAAAA9555552AAAAD5555AAAA5555AAA9555AAAD552AAD55AAB552AB552A954AA552A956A956A952AD5AB56AD5AB52A56AD4AD4AD4AD6A56B5294AD6B5AD6B5AD6B4A52D6B4A5A52D29696B4B4B4B4B4B69696D2DA5B49692DB496DA496DA4925B6DB6D24924924DB6DB";
defparam ram_block1a77.mem_init2 = "6C924DB64936C936C9B64D9364D9364D9B264C993264C99B32664CC999B333366666666CCCCCCE666666673333999CCC6673398CC67318CE7318C6318C631CE718E718E31C718E38E38E38E38E3C71E38F1E3870E1E3C38787870F878787C3C1E0F87C1F07C1F03E07C0FC0FE07F03FC07F00FF807FC00FFC003FFC000FFFF000007FFFFFFFE000000000001FFFFFFFF800007FFF8001FFE003FF007FC03FC03F80FE03F03F03E07C0F83E0F87C1E1F0F0787878F0F1E1C3870E3C70E38E38E38E38E31C738C738C6318C6319CC673198CC667333399999999999999B333666CCD9B366CD9326C9B24D926D9249B6DB6DB6DB6D24B6D25B49692D2D2D2D2D694";
defparam ram_block1a77.mem_init1 = "B5AD6B5AD6A56B52A56AD5AA55AA552AB556AA95552AAAAD555555555555555555556AAAAD555AAA554AAD56A956AD5AB52B52B5294A5294B5A52D2D2D2D2DA5B492DB492496DB64924DB649B64D9364C9B3264CD99933332666666733331998CC67319CE6318E738C738E39C71C78E3871E3C78F0F1E1F0F0F87C1F07C1F81F81F80FE01FF007FE003FFF80000FFFFFFFFFFFFFFFFFC00007FFE001FF803FC03F80FC0FC0F81F0783E1E0F0F0F1E1C3870E3871C71C738E31CE318C6339CC66331999CCCCCCCCCCD99933264C99326C9B649B6492492492496DA4B69692D29696B5A5295AD4AD4AD5AA55AAD54AA95552AAAAB555555555556AAAAA5556AAD5";
defparam ram_block1a77.mem_init0 = "4AA55AB56AD4AD6A5294A5AD2D2D2D2DA4B692496DB6D9249B64DB26CD9B366CCD9999999999999CCC663398C6318C738E71C71C71E3870E1C3C3C3C1E0F07C0F81F81FC07F803FE001FFFC0000003FFFFE0000001FFFC007FE00FF01FC0FC0F83E0F8783C3C3C78F1E3871C71C738E718C6319CE67339999CCCCCD999933264C993649B24DB6DB6DB6DA4B692D2D2D2D694A52B5A95AB56A954AAD552AAAB55555555555554AAAAD552AB55AB54AD4AD4A5294B5A5A5A5A4B6924B6DB6C924DB26C9B366CC999B33333333999CCE6339CE738C71CE38E3C70E3C3878787C3E0F83F03F01FC03FE003FFE000003FFFFFFE000003FFE003FE01FC07E07C0F87C1";

cyclonev_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 8191;
defparam ram_block1a5.port_a_logical_ram_depth = 65536;
defparam ram_block1a5.port_a_logical_ram_width = 24;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init3 = "07C3E07C0FC07F00FF800FFF800000FFFFFFF800000FFF800FF807F01F81F83E0F87C3C3C3878E1C78E38E71C639CE7398CE6733399999999B33266CD9B26C9B64926DB6DA492DA4B4B4B4B5A5294A56A56A55AB55AA9556AAAA55555555555555AAAA9556AA552AD5AB52B5A94A52D696969692DA4B6DB6DB6DB649B24D93264C9993333666667333399CCE7318C631CE39C71C71C38F1E3C7878783C3E0F83E07E07F01FE00FFC007FFF0000000FFFFF80000007FFF000FF803FC07F03F03E07C1E0F078787870E1C38F1C71C71CE39C6318C63398CC6673333333333333666CD9B366C9B64DB24936DB6D2492DA4B696969696B4A5294AD6A56AD5AB54AA5";
defparam ram_block1a5.mem_init2 = "56AAD554AAAAAD55555555555AAAAA95552AA556AB54AB56A56A56B5294B5AD2D29692D2DA4B6D24924924924DB24DB26C993264C99933366666666667333198CC67398C6318E718E39C71C71C38E1C3870F1E1E1E0F0F83C1F03E07E07E03F807F803FF000FFFC00007FFFFFFFFFFFFFFFFE00003FFF800FFC01FF00FE03F03F03F07C1F07C3E1E1F0F1E1E3C78F1C38E3C71C738E39C639CE318CE7319CC6633319999CCCCCCC99999333664C99B264D9364DB24DB64924DB6D24925B6925B4B69696969694B5A5294A5295A95A95AB56AD52AD56AA554AAB5556AAAAD555555555555555555556AAAA95552AAD55AA954AB54AB56AD4A95AD4AD6B5AD6B5A";
defparam ram_block1a5.mem_init1 = "52D69696969692D25B496DA496DB6DB6DB6DB24936C93649B26C99366CD9B3666CCD999B333333333333339999CCC663319CC67318C6318C639C639C718E38E38E38E38E1C78E1C3870F1E1E3C3C3C1E1F0F07C3E0F83E07C0F81F81F80FE03F807F807FC01FF800FFF0003FFFC00003FFFFFFFF000000000000FFFFFFFFC00001FFFE0007FF8007FE007FC03FE01FC07F81FC0FE07E07C0F81F07C1F07C3E0F0787C3C3C3E1C3C3C3878F0E1C38F1E38F1C78E38E38E38E38E31C718E31CE31CE718C6318C6319CE6319CC663399CCC6673339999CCCCCCCCE666666CCCCCCCD9999B332664CC99B3264C993264C9B364D9364D9364DB26D926D924DB64926D";
defparam ram_block1a5.mem_init0 = "B6DB6492492496DB6DB4924B6D24B6D25B692D25B4B696D2D2DA5A5A5A5A5AD2D29694B4A5AD694A5AD6B5AD6B5AD6A5295AD4AD6A56A56A56AD4A95AB56AD5AB56A952AD52AD52A954AA552A955AA955AAB556AA9556AAB5552AAB5554AAAB55556AAAA9555552AAAAAAD555555554AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA95555555556AAAAAAA5555556AAAAAD55556AAAAD5554AAAA5555AAAB5556AAAD554AAA5552AA9556AA9556AA9552AA554AA9552AB556AA556AA556AB552AB55AAD54AA552A954AA55AAD56A954AA55AA552AD52A956A956A956A956A956A956A956AD52AD52AD5AA55AB54AB56A952AD52A55AB54A956AD52AD5AA";

cyclonev_ram_block ram_block1a29(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.clk0_output_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "rom";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "clock0";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 8192;
defparam ram_block1a29.port_a_first_bit_number = 5;
defparam ram_block1a29.port_a_last_address = 16383;
defparam ram_block1a29.port_a_logical_ram_depth = 65536;
defparam ram_block1a29.port_a_logical_ram_width = 24;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init3 = "FFFFFFF000FF807F03F07C1E1E1E1C38E1C738E739CE63319999999933264D936C924924B6D2D2D2D6B5AD4AD52AD54AAA95555555554AAA955AAD5A95A94A5A52DA5B49249249364993664CCCD9CCCCC67318C639C71C71C387878783E0F81FC07F800FFFE0000000003FFF800FF01FC0F83E0F0F0F1E3C71C71CE318C673399999999993264D936492492496D25A5AD294A56A54AB552AA95555555555552AA955AA54AD4A5296B4B496D24924924DB264D993332666333198CE738C738E3871E3C3C3C3E0F81F80FE00FFF00000FFFFF800003FF803FC0FC0F83E1F0F1E1C38E38E39C6319CC6633333333666CD9364DB24924B6D25A5A5AD295A95AB54AA";
defparam ram_block1a29.mem_init2 = "555AAAAAAAAAAAAAAD552A956AD4AD4A5AD2D2D25B4924926D926CD93366666666663319CE738C71C71C78F0E1E0F07C1F81F807FC007FFFC00000003FFFE003FE03F81F83E0F0F0F0E1C38E38E71CE7398CC6666666666CC99364D924DB6D24B692D2D694A52B52A55AAD552AAAAB5555AAAAA9556AB54A95A94A52D69692D24B6DB6C926C9B366CCD9999998CCE6339CE31C638F1C78F0E0F0F87C0FC0FE01FF000FFFFFE0003FFFFF8007FC03F81F83E0F8787878F1C78E31C639CE63399CCCCCCCCC99B366C936C924924B6D2DA5AD294A52B52AD52A9554AAAAAAAAAAAAAA5552A956AD5A94A5296B4B696D24924924DB26C99336664CCCC6663319CE73";
defparam ram_block1a29.mem_init1 = "8C71C71C70E1C3C3C1E0F83F03F807FC007FFFC000000007FFFC003FE03F81F81F0787C3C7870E38E38E31CE7398CE667333333666CC9B3649B6C92492DB4B69696B4A52B52B56A954AAB55556AAAAAAB55556AA954AB56AD6A5294B4B4B496D24924924DB26C9932666CCCCCCE667319CE738C718E3C71E3C78787C3E0F81F80FE00FFC001FFFFFFFFFFFFFE0007FE00FE03F07E0F87C3C3C78F1C38E38C738C6319CCE66633336666CC99326D936DB6DB6DA4B6969696B5AD6A56AD5AAD54AAA555555555555555AAAD54AA54A95A94A52D6969692DA496DB64926C9326CD993333333333399CCE739CE31C71C71C38F0E1E1F0F83E0FC0FE03FC00FFF8000";
defparam ram_block1a29.mem_init0 = "00FFFFF000001FFF003FC07F03F07E1F0787878F1E3871C718E31CE7319CC6667333332666CC99364D926DB6DB6DB496D2D2D2D6B4AD6A56AD5AA556AA955554AAAAAAA955556AA955AA55AB52B5AD6B4A5A5A5B496DB6DB6DB649B26CD9B36666CCCCCC6663319CC631CE31C71C71C38F0E1E1E0F0781F03F03F807FC007FFE000000000000000FFFE007FC03F80FC1F83E0F0F878F0E1C38E38E38E718E7318CE673339999999333664C993649B64926DA4925B496969696B5AD6B52B52AD5AAD55AAA9555555AAAA5555556AAA554AA55AB52B52B5AD296B4B4B696DA492DB64926D926CD93266CCD999999999CCC66339CE739C638E31E38E1C78F0F0F0F";

cyclonev_ram_block ram_block1a102(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a102_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a102.clk0_core_clock_enable = "ena0";
defparam ram_block1a102.clk0_input_clock_enable = "ena0";
defparam ram_block1a102.clk0_output_clock_enable = "ena0";
defparam ram_block1a102.data_interleave_offset_in_bits = 1;
defparam ram_block1a102.data_interleave_width_in_bits = 1;
defparam ram_block1a102.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a102.init_file_layout = "port_a";
defparam ram_block1a102.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a102.operation_mode = "rom";
defparam ram_block1a102.port_a_address_clear = "none";
defparam ram_block1a102.port_a_address_width = 13;
defparam ram_block1a102.port_a_data_out_clear = "none";
defparam ram_block1a102.port_a_data_out_clock = "clock0";
defparam ram_block1a102.port_a_data_width = 1;
defparam ram_block1a102.port_a_first_address = 32768;
defparam ram_block1a102.port_a_first_bit_number = 6;
defparam ram_block1a102.port_a_last_address = 40959;
defparam ram_block1a102.port_a_logical_ram_depth = 65536;
defparam ram_block1a102.port_a_logical_ram_width = 24;
defparam ram_block1a102.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a102.ram_block_type = "auto";
defparam ram_block1a102.mem_init3 = "D56AA556AA9555AAAAD555556AAAAAAAAAAAAAAAAAB555555AAAAD554AAB556AA552A956AD52A54AD5A95AD4AD6B5AD6B5A52D696B4B4B4B49696D25B496DA4925B6DB6DB6DB24936D926D936C9B26CD93264C9933666CCD9999333333333333339999CCCE663319CC67318C6739C6318E718E71C638E38E38E38E3871C3871E3C7870F0F1E1E1F0F0F87C3E0F07C1F83E07C0FC0FE07F01FC07F807FC01FF800FFE000FFFE00003FFFFFF0000000000000000000FFFFFFE00003FFF8003FFC007FE00FF807F80FF01FC0FE07E07E0FC1F03E0F87C1F0F8783C3C3C3C3C3C3878F1E3C78E1C78E3871C71C71C718E38C718E718E739C6318CE7398CE63398CC6";
defparam ram_block1a102.mem_init2 = "67331999CCCCCE66666666666CCCCCD999333664CD993264C9B364D9B26D93649B649B64936DB6C924924924B6DB6924B6925B496D2DA5A4B4B4B4B4B5A5AD2D6B4A52D6B5A94A52B5295A95A952B56AD5AA54AB54AA552AB552AB554AAB5552AAAD55552AAAAA9555555555555555555555555556AAAAAA55554AAAB5552AA9556AAD54AAD56AB54AB54AB56AD5AB56A56AD4AD6A56B5294A5294A5294B5AD2D694B4B4A5A5A5B4B4B49692D25B496DA4B6D2496DB6D24924924924936DB64926DB24DB24DB26C9364D9366C9B364C993264C99B3266CCD999333266664CCCCCCCCCCCCCCCCCCCCE66663333999CCC6673398CC67319CC6339CC6318C6318C6";
defparam ram_block1a102.mem_init1 = "31CE718E718E71CE38C71C638E38E38E38E38E3871C70E3871E3870E1C3870E1E3C387870F0F0F0F0F0F0F8787C3C1E0F07C3E0F87C1F07C0F83E07C0F81F81F81F81F80FC07E03F80FF01FE03FC01FE00FF803FE007FE003FF8007FFC001FFF80007FFFC00003FFFFF80000003FFFFFFFFFFFFFC00000000003FFFFFFFFFFFFFC00000007FFFFF00000FFFFC0003FFF8001FFF0007FF000FFE007FE007FC00FF807FC03FC03FC03FC07F01FE07F01FC0FE07F03F03F03F03F03E07C0F81F03E0F81F07C1F07C1E0F83C1F0F83C1E0F0787C3C1E1E0F0F0F0F0F87870F0F0F0F1E1E1C3C7878F1E1C3878F1E3C78F1C3871E3871E3871C38E1C71C38E38F1C71";
defparam ram_block1a102.mem_init0 = "C71C70E38E38C71C71C71C638E38C71C638E71C638C718E31CE39C639C639CE31CE718C639CE718C6318C6318C6318C6339CE7318C67398C67318CE63398CE63398CE67319CCE673198CC6633199CCE66333998CCE667333999CCCC6667333399998CCCCC6666673333331999999999CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC9999999999B33333326666664CCCCC99999B333366664CCCD999933326664CCC999B3336664CC999B332664CC999B33666CCD99332664CD99B33664CD99B3266CC99B3266CCD9B3266CC99B3266CD9933664C99B3664CD9B3264CD9B3264CD9B3264C99B3664C993366CD993264CD9B366CC993266CD9B3664C9932";

cyclonev_ram_block ram_block1a126(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a126_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a126.clk0_core_clock_enable = "ena0";
defparam ram_block1a126.clk0_input_clock_enable = "ena0";
defparam ram_block1a126.clk0_output_clock_enable = "ena0";
defparam ram_block1a126.data_interleave_offset_in_bits = 1;
defparam ram_block1a126.data_interleave_width_in_bits = 1;
defparam ram_block1a126.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a126.init_file_layout = "port_a";
defparam ram_block1a126.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a126.operation_mode = "rom";
defparam ram_block1a126.port_a_address_clear = "none";
defparam ram_block1a126.port_a_address_width = 13;
defparam ram_block1a126.port_a_data_out_clear = "none";
defparam ram_block1a126.port_a_data_out_clock = "clock0";
defparam ram_block1a126.port_a_data_width = 1;
defparam ram_block1a126.port_a_first_address = 40960;
defparam ram_block1a126.port_a_first_bit_number = 6;
defparam ram_block1a126.port_a_last_address = 49151;
defparam ram_block1a126.port_a_logical_ram_depth = 65536;
defparam ram_block1a126.port_a_logical_ram_width = 24;
defparam ram_block1a126.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a126.ram_block_type = "auto";
defparam ram_block1a126.mem_init3 = "0000000000FFFF8003FF803FE01FE03F03F83F07C1F07C3E1E1E1E1E3C78F1E38E1C71C738E31CE318C6318CE633198CCCC6666666666CCCD993366CD9366D936C936D92492492DB6925B49696969696B4A5AD6B5295A95AB56AD52AD54AAD556AAA9555555AAAAAAAAAD555554AAAB554AA955AA55AB56AD4AD4A56B5AD296B4B4B4B4B696D24B6DA4924924DB6493649B26CD9B366CC99993333333333339998CC67319CC6318E738C71CE38E38E3C70E3C78F0F0E1F0F0F87C1F07C0F81F80FE03FC03FE007FF8000FFFFF0000000000000007FFFFC000FFF003FE00FE01F80FC0FC1F03E1F0787C3C3C3C7870E1C78E3871C738E39C639CE739CE63398CC";
defparam ram_block1a126.mem_init2 = "666333333333333336664CD9B366C9B26C9B649B6DB24924B6DB496D25B4B4B4B4B4A5AD6B5AD4A56A56AD5AB55AA556AAD552AAA95555554AAAAAAAD5555556AAA9554AA955AA55AA54A95A95AD4A5294A5AD2D2D2D2D25A4B6D24B6DB6DB6D924DB64DB26C99366CC99B336666664CCE66666733198CC67398C631CE718E39C71C71C70E3870E1C3C7878783C3E1F07C1F03F07F03F80FF00FF801FFC001FFFF0000000007FE0000000007FFFC001FFC00FF807F80FE07F07E07C1F07C3E1F0F0F0F0E1E3C78E1C70E38E38C71CE39CE318C63398CE6333999CCCCCCCCCCCCCD99933264C99326C9B24D924DB6C92492496DB492DA5B4B49694B4B5A5294A5";
defparam ram_block1a126.mem_init1 = "295A95A95AB56A956AB552AA5552AAA95555554AAAAAAAA55555552AAA9554AA955AAD56AD52B56A56A56B5AD6B5A52D2969696D2DA4B6925B6DA4924DB6D924DB26C9326C993264CD99933332666666733331998CC67319CE6318E738C738E31C71C71C38E1C78F0E1E3C3C3C1E1F0F83E0F83F03E03F01FC07F803FE003FF8001FFFFC000000000000000000007FFFE0007FF800FF803FC07F01FC0FC1F83F07C3E0F078783C387870F1E3871E38E38E38E38C718E718C6318C67319CCE67333199999999999999333666CD99366C993649B24DB24936DB6DB6DA492DB496D2DA5A5A5A5A52D694A5294AD6A56A56AD5AA54AA552AB556AAB5554AAAAAD555";
defparam ram_block1a126.mem_init0 = "5555555555554AAAAAD5552AA9552AB55AAD52A54A952B52B5A94A5294B5A52D2969692D2DA5B692DB4924924924924DB649B64D9364D93264C99B32666CCCCC9999999CCCCCE6673399CC67318C6318C639C638C71C71C71C71C38E1C3870E1E1C3C3C1E1E0F07C3E0FC1F03F03F03F80FE01FE00FFC00FFF0007FFFC000001FFFFFFFFFFFFFFF0000007FFFC000FFE003FE00FF80FF01F80FC0FC0F81F07C1F0F87C3C1E1E1E1C3C7870E3C78E3871C71C71C638E718E718C6318C63398CE633199CCCE66666673366666664CCC99B3266CD9B264D9364DB26D924DB6C924924924B6DA496DA4B49692D2D2D2D29694B5AD6B5AD6B52B52B52B56AD5AA55AA";

cyclonev_ram_block ram_block1a150(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a150_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a150.clk0_core_clock_enable = "ena0";
defparam ram_block1a150.clk0_input_clock_enable = "ena0";
defparam ram_block1a150.clk0_output_clock_enable = "ena0";
defparam ram_block1a150.data_interleave_offset_in_bits = 1;
defparam ram_block1a150.data_interleave_width_in_bits = 1;
defparam ram_block1a150.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a150.init_file_layout = "port_a";
defparam ram_block1a150.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a150.operation_mode = "rom";
defparam ram_block1a150.port_a_address_clear = "none";
defparam ram_block1a150.port_a_address_width = 13;
defparam ram_block1a150.port_a_data_out_clear = "none";
defparam ram_block1a150.port_a_data_out_clock = "clock0";
defparam ram_block1a150.port_a_data_width = 1;
defparam ram_block1a150.port_a_first_address = 49152;
defparam ram_block1a150.port_a_first_bit_number = 6;
defparam ram_block1a150.port_a_last_address = 57343;
defparam ram_block1a150.port_a_logical_ram_depth = 65536;
defparam ram_block1a150.port_a_logical_ram_width = 24;
defparam ram_block1a150.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a150.ram_block_type = "auto";
defparam ram_block1a150.mem_init3 = "AB54AB56AD5A95A95A95AD6B5AD6B5A52D29696969692D25A4B6D24B6DA4924924926DB64936C9B64D9364C9B366CC99B326664CCCCCCD99CCCCCCCE66733198CE63398C6318C631CE31CE38C71C71C71C38E3C78E1C3C7870F0F0F0787C3E1F07C1F03E07E07E03F01FE03FE00FF800FFE0007FFFC000001FFFFFFFFFFFFFFF0000007FFFC001FFE007FE00FF00FE03F81F81F81F07E0F87C1E0F0F0787870F0E1C3870E3871C71C71C71C638C738C6318C6319CC673399CCCE66667333333266666CCC99B3264C99364D9364DB24DB64924924924925B692DB4B69692D2D29694B5A5294A52B5A95A952A54A956AB55AA9552AA95556AAAAA5555555555555";
defparam ram_block1a150.mem_init2 = "5556AAAAA5555AAAD55AA954AA54AB56AD4AD4AD6A5294A52D694B4B4B4B4B696D25B6924B6DB6DB6D9249B649B24D9326CD93366CCD999333333333333331999CCE67319CC6318C631CE31C638E38E38E38F1C38F1E1C3C38783C3C1E0F87C1F83F07E07F01FC07F803FE003FFC000FFFFC000000000000000000007FFFF0003FF800FF803FC07F01F80F81F83E0F83E1F0F0787878F0E1E3C70E3871C71C718E39C639CE318CE7319CC6633319999CCCCCCC99999333664C99326C9926C9B64936DB64924B6DB492DA4B696D2D2D29694B5AD6B5AD4AD4AD5A956AD56AB552AA5552AAA95555554AAAAAAAA55555552AAA9554AA955AAD52AD5AB52B52B529";
defparam ram_block1a150.mem_init1 = "4A5294B5A5A52D25A5B4B6925B6D24924926DB6493649B26C993264C99933366666666666667333998CE63398C6318E738E71C638E38E1C70E3C78F0E1E1E1E1F0F87C1F07C0FC1FC0FE03FC03FE007FF0007FFFC000000000FFC000000001FFFF0007FF003FE01FE03F81FC1F81F07C1F0F8783C3C3C7870E1C38E1C71C71C738E31CE718C6339CC6633199CCCCCCE664CCCCCD99B3266CD9326C9B64DB64936DB6DB6DA496DA4B49696969696B4A5294A56B52B52A54AB54AB552AA5552AAAD5555556AAAAAAA55555552AAA9556AAD54AB55AB56AD4AD4A56B5AD6B4A5A5A5A5A5B496D25B6DA49249B6DB24DB26C9B26CD9B3664CCD99999999999998CCC";
defparam ram_block1a150.mem_init0 = "663398CE739CE738C738E39C71C38E3C70E1C3C7878787C3C1F0F81F07E07E03F00FE00FF801FFE0007FFFFC000000000000001FFFFE0003FFC00FF807F80FE03F03E07C1F07C3E1E1F0E1E1E3C78E1C78E38E38E71C639CE318C67319CC663333999999999999333266CD9B366C9B24D924DB64924924B6DA496D2DA5A5A5A5AD296B5AD4A56A56AD5AB54AB552AA555AAAA5555556AAAAAAAAB5555552AAAD556AA556A956AD5AB52B5295AD6B4A5AD2D2D2D2D25B492DB6924924936D926D936CD9366CD99336666CCCCCCCCCC666633198CE6318C6318E718E39C71C70E38F1E3C78F0F0F0F0F87C1F07C1F83F81F80FF00FF803FF8003FFFE0000000000";

cyclonev_ram_block ram_block1a174(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a174_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a174.clk0_core_clock_enable = "ena0";
defparam ram_block1a174.clk0_input_clock_enable = "ena0";
defparam ram_block1a174.clk0_output_clock_enable = "ena0";
defparam ram_block1a174.data_interleave_offset_in_bits = 1;
defparam ram_block1a174.data_interleave_width_in_bits = 1;
defparam ram_block1a174.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a174.init_file_layout = "port_a";
defparam ram_block1a174.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a174.operation_mode = "rom";
defparam ram_block1a174.port_a_address_clear = "none";
defparam ram_block1a174.port_a_address_width = 13;
defparam ram_block1a174.port_a_data_out_clear = "none";
defparam ram_block1a174.port_a_data_out_clock = "clock0";
defparam ram_block1a174.port_a_data_width = 1;
defparam ram_block1a174.port_a_first_address = 57344;
defparam ram_block1a174.port_a_first_bit_number = 6;
defparam ram_block1a174.port_a_last_address = 65535;
defparam ram_block1a174.port_a_logical_ram_depth = 65536;
defparam ram_block1a174.port_a_logical_ram_width = 24;
defparam ram_block1a174.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a174.ram_block_type = "auto";
defparam ram_block1a174.mem_init3 = "993264CD9B366CC993266CD9B3664C993366CD993264CD9B3264C99B3664C99B3664C99B3664CD9B3264CD993366CC99B3266CC99B3666CC99B3266CC99B33664CD99B33664CC99933666CCD99B332664CC999B332664CCD999B3326664CCC9999333366664CCCD9999B33332666664CCCCCC9999999B33333333326666666666666666666666666666666666666666673333333331999999CCCCCC66666333339999CCCC6667333999CCCE66333998CCE6733198CC663319CCE67319CCE63398CE63398CE6319CC6339CC6319CE7398C6318C6318C6318C631CE738C631CE718E738C738C738E718E31C638C71CE38C71C638E38C71C71C71C638E38E1C71C7";
defparam ram_block1a174.mem_init2 = "1C71E38E3871C70E3871C38F1C38F1C3871E3C78F1E3C3870F1E3C3C7870F0F1E1E1E1E1C3C3E1E1E1E1E0F0F0787C3C1E0F0783E1F0783E0F07C1F07C1F03E0F81F03E07C0F81F81F81F81F81FC0FE07F01FC0FF01FC07F807F807F807FC03FE007FC00FFC00FFE001FFC001FFF0003FFF80007FFFE00001FFFFFC00000007FFFFFFFFFFFFF800000000007FFFFFFFFFFFFF80000003FFFFF800007FFFC0003FFF0007FFC003FF800FFC00FF803FE00FF007F80FF01FE03F80FC07E03F03F03F03F03E07C0F83E07C1F07C3E0F87C1E0F0787C3C3E1E1E1E1E1E1E1C3C3878F0E1C3870E1C38F1C38E1C71C38E38E38E38E38E38C71C638E71CE31CE31CE718";
defparam ram_block1a174.mem_init1 = "C6318C6318C67398C67319CC663399CCC6673339998CCCCE666666666666666666664CCCC9999333666CC99B3264C993264D9B26CD9364D926C9B649B649B6C924DB6D92492492492496DB6D2496DA4B6D25B49692D25A5A5B4B4B4A5A5A52D696B5A5294A5294A5295AD4AD6A56AD4AD5AB56AD5AA55AA55AAD56AA556AAD552AA9555AAAA55554AAAAAAD555555555555555555555555552AAAAA955556AAA9555AAA555AA955AA954AA55AA54AB56AD5A952B52B5295A94A52B5AD694A5AD696B4B5A5A5A5A5A4B4B696D25B492DA492DB6DA4924924926DB6D924DB24DB24D936C9B364D9B264C9933664CD999333666666CCCCCCCCCCCE66667333199CC";
defparam ram_block1a174.mem_init0 = "C663398CE6339CE6318C739CE31CE31C638E31C71C71C71C38E3C70E3C78F1E3C387878787878783C3E1F07C3E0F81F07E0FC0FC0FE07F01FE03FC03FE00FFC007FF8003FFF80000FFFFFFE0000000000000000001FFFFFF80000FFFE000FFE003FF007FC03FC07F01FC0FE07E07C0F83F07C1E0F87C3E1E1F0F0F1E1E1C3C78F1C3871C38E38E38E38E38C71CE31CE318C739CC6319CC673198CCE6673333999999999999993333666CCD993264C99366C9B26D936C936D9249B6DB6DB6DB4924B6D25B496D2D25A5A5A5AD2D694B5AD6B5AD6A56B52B56A54A956AD52A954AAD55AAA5556AAAB555555AAAAAAAAAAAAAAAAAAD555556AAAB5552AAD54AAD56";

cyclonev_ram_block ram_block1a54(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a54_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a54.clk0_core_clock_enable = "ena0";
defparam ram_block1a54.clk0_input_clock_enable = "ena0";
defparam ram_block1a54.clk0_output_clock_enable = "ena0";
defparam ram_block1a54.data_interleave_offset_in_bits = 1;
defparam ram_block1a54.data_interleave_width_in_bits = 1;
defparam ram_block1a54.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a54.init_file_layout = "port_a";
defparam ram_block1a54.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a54.operation_mode = "rom";
defparam ram_block1a54.port_a_address_clear = "none";
defparam ram_block1a54.port_a_address_width = 13;
defparam ram_block1a54.port_a_data_out_clear = "none";
defparam ram_block1a54.port_a_data_out_clock = "clock0";
defparam ram_block1a54.port_a_data_width = 1;
defparam ram_block1a54.port_a_first_address = 16384;
defparam ram_block1a54.port_a_first_bit_number = 6;
defparam ram_block1a54.port_a_last_address = 24575;
defparam ram_block1a54.port_a_logical_ram_depth = 65536;
defparam ram_block1a54.port_a_logical_ram_width = 24;
defparam ram_block1a54.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a54.ram_block_type = "auto";
defparam ram_block1a54.mem_init3 = "54AB54A952A56A54A56A5294A5294A5AD2D696969696D2DA5B492DA4925B6DB6DB6D9249B6C93649B26C9B364C993266CCD999B33333266673333331998CCE673198C6739CE739CE31CE31C738E38E38E3C71C38F1E3C3878F0F0F0F8783C1E0F83E0FC1F81F81F80FE01FC01FE007FF001FFF80003FFFFFE000000000000000FFFFFF80003FFE001FFC01FF00FF01FC07E07E07E0F81F0783E1F0F0787878F0F1E3C78F1C38E38E38E38E39C738C739CE739CE63398CC6633319999CCCCCCCC99999B33666CD9B366C9B36C9B24DB249B6DB6DB6DB6DA496DA4B49692D2D2D69694A5AD6B5AD4A56A56AD5AB56A956AA556AAD556AAAD55555AAAAAAAAAAAAA";
defparam ram_block1a54.mem_init2 = "AAA9555552AAA5552AA556AB55AA54A952B52B52B5AD6B5AD296B4B4B4B4B4B692DA4B6DA4924924926DB649B64DB26C99366CD99332666CCCCCCCCCCCCCCC66633198CE6339CE739CE31CE39C71C71C71C70E3870E1E3C3C78783C3E1F0F83E07C1F81F80FE03F807FC01FFC007FFE00003FFFFFFFFFFFFFFFFFFFF80000FFFC003FF007FC03F80FE07F03E07C1F07C1E0F0F8787870F0E1C38F1C78E38E38E71C639C639CE7318CE63399CCCE6666333333366666CCC99B366CD9326C93649B6C924DB6DB492496D24B49692D2D2D696B4A5294A52B52B52B56A952A956AA555AAAD5552AAAAAA9555555552AAAAAAD5556AAB556AA552AD52A54AD4AD4AD6";
defparam ram_block1a54.mem_init1 = "B5AD6B4A5A52D2D25A4B496DA492DB6DB6DB249B6C9B64D9366CD9B3664CCD99999999999999CCCE673198C6739CE718C718E39C71C71E38E1C3870E1E1E1E1E0F0783E0F83F07E03F01FC03FC01FF800FFF80003FFFFFFFF8000FFFFFFFFE0000FFF8007FC01FF01FC07E03F07E0F83E0F0783C3C3C3878F1E3C70E38E38E38E71CE318E739CC63399CCE663333339999333332664CD99326CD93649B24DB6C924924925B6925B4B69696969694B5AD6B5A94AD4AD5AB54AB54AAD55AAAD5552AAAAAAD55555552AAAAAAD5556AA9552AB55AA54A952B52B5294A5294B5A5A5A5A5A4B492DA4925B6DB6C924DB24D926CD93264C99B33266666666666667333";
defparam ram_block1a54.mem_init0 = "99CC67318CE718C738C71C638E3871C38F1E3C387878787C3E0F07C0F81F81F80FF01FF007FE001FFF800007FFFFFFFFFFFFFFE00000FFFC003FF007F807F01FC0FC1F83E0F83C1E1F0F0E1E1C3870E3871C71C718E39C631CE7398C673399CCCE6666666666664CCD993366C99364DB26D9249B6DB6DB6925B692DA5A5A5A5A52D694A52B5A95A952A54AB54AAD54AAA5554AAAAAAD555555555AAAAAA95552AA955AA956A956AD4AD4AD6A5294B5AD2D2D6D2D2DA4B6924B6DB6DB6C926DB26D9366C993266CC999933333333331999CCE67319CE739CE718E71C638E38E1C70E3C7870F0F0F0F0783E0F83E07C0FE07F00FF00FFC007FFC0001FFFFFFFFFF";

cyclonev_ram_block ram_block1a78(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a78_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a78.clk0_core_clock_enable = "ena0";
defparam ram_block1a78.clk0_input_clock_enable = "ena0";
defparam ram_block1a78.clk0_output_clock_enable = "ena0";
defparam ram_block1a78.data_interleave_offset_in_bits = 1;
defparam ram_block1a78.data_interleave_width_in_bits = 1;
defparam ram_block1a78.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a78.init_file_layout = "port_a";
defparam ram_block1a78.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a78.operation_mode = "rom";
defparam ram_block1a78.port_a_address_clear = "none";
defparam ram_block1a78.port_a_address_width = 13;
defparam ram_block1a78.port_a_data_out_clear = "none";
defparam ram_block1a78.port_a_data_out_clock = "clock0";
defparam ram_block1a78.port_a_data_width = 1;
defparam ram_block1a78.port_a_first_address = 24576;
defparam ram_block1a78.port_a_first_bit_number = 6;
defparam ram_block1a78.port_a_last_address = 32767;
defparam ram_block1a78.port_a_logical_ram_depth = 65536;
defparam ram_block1a78.port_a_logical_ram_width = 24;
defparam ram_block1a78.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a78.ram_block_type = "auto";
defparam ram_block1a78.mem_init3 = "66CD9B3264C993366CD9B3264C99B366CC993266CD9B3264CD9B3664C99B3664C99B3664C99B3664CD9B3266CD9933664CD993266CC99B3266CCD9933664CC99B32664CD99B33664CC999332664CC999B336664CC999B332666CCCD999B3336666CCCD99993333266664CCCCD99999B33333266666664CCCCCCCCC9999999999999999999999999999999999999999999CCCCCCCCCE66666673333319999CCCCC666633339998CCC666333199CCC66733198CCE673399CCE673198CE67319CC67319CC67319CE6339CC6339CE6318CE739CE739CE739CE739CE318C639CE318E718C738C738C718E71CE39C738E71C738E39C71C638E38E38E31C71C71C38E38";
defparam ram_block1a78.mem_init2 = "E38E3C71C70E38F1C78E3C70E3C70E3C78E1C3870E1C3878F1E1C3C7878F0F0E1E1E1E1C3C3C3E1E1E1E1F0F0F8783C3E1F0F87C3E0F07C1F0F83E0F83E0FC1F07E0F81F03F07E07E07E07E07E03F01F80FE07F01FE03F807F80FF807F803FC01FF803FF003FF001FFC003FFE000FFFC000FFFF80003FFFFC000003FFFFFFF00000000000001FFFFFFFFFFFE00000000000007FFFFFFE000003FFFF80003FFFC000FFFC003FFC007FF003FF007FE01FF007F807F00FE01FC07F03F80FC0FC0FC0FC0FC1F83F07C0F83E0F83E1F0783E1F0F8783C3C1E1E1E1E1E1E1E3C3C7870F1E3C78F1E3C70E3C71E38E1C71C71C71C71C71C738E39C718E31CE31CE318E7";
defparam ram_block1a78.mem_init1 = "39CE739CE7398C63398CE63399CC66333998CCE66633333199999999999999999999B33336666CCC99933664CD9B366CD9B264D9B26C9B26D93649B649B64936D924926DB6DB6DB6DB692492DB6925B692DA4B696D2DA5A5B4B4B4B5A5A5AD2D694A5AD6B4A52B5AD6A52B5295A952B52A54A952A55AB55AA552A955AA9552AAD552AAB5555AAAAB5555552AAAAAAAAAAAAAAAAAAAAAAAAAAD555554AAAA95556AAA555AAA554AAD56AB55AA55AB54A952A56AD4AD4AD6A56B5A94A5296B5AD296B4B4A5A5A5A5A5B4B49692DA4B6925B6D2492DB6DB6DB6DB24926DB249B64DB26C9364C9B264D9B366CC99B32664CCC99999933333333333199999CCCE6633";
defparam ram_block1a78.mem_init0 = "399CC67319CC6319CE739C631CE31CE39C718E38E38E38E3871C38E1C3870E1C3C7878787878787C3C1E0F87C1F07C0F81F03F03F01F80FE03FC03FC01FF003FF8007FFC0007FFFE0000003FFFFFFFFFFFFFFFFFFE0000007FFFF0001FFF000FFC00FF803FC03F80FE03F81F81F83F07E0F83E1F0783C1E1E0F0F0E1E1E3C3870E1C78E3C71C71C71C71C738E31CE31CE718C6339CE63398CE6733199CCCCC66666666666666CCCC999B3266CD99366C99364D926C936C936DB2492492492496DB492DA4B692D2DA5A5A5A52D296B4A5294A5295A94AD4A95AB56AD52AD56AB552AA555AAA95554AAAAAB5555555555555555556AAAAA95554AAAD552AA552AB";

cyclonev_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 8191;
defparam ram_block1a6.port_a_logical_ram_depth = 65536;
defparam ram_block1a6.port_a_logical_ram_width = 24;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init3 = "AA954AA9556AAA55552AAAAAD555555555555555555AAAAAA55552AAB554AA955AAD56A956AD5AB52A56A52B5294A5294A5AD29694B4B4B4B69692DA4B6925B6D249249249249B6D926D926C9364D9326CD93366CC99B3326666CCCCCCCCCCCCCC6666733199CCE63398CE7398C631CE718E718E39C71C71C71C71C78E3C70E1C3878F0F0E1E1E0F0F0783C1F0F83E0FC1F83F03F03F80FE03F807F803FE007FE001FFF0001FFFFC000000FFFFFFFFFFFFFFFFFFF8000000FFFFC0007FFC003FF801FF007F807F80FE03F01F81F81F03E07C1F07C3E0F0787C3C3C3C3C3C3C7870E1C3870E3871C38E38E38E38E31C738E718E718C739CE7318C67319CC67339";
defparam ram_block1a6.mem_init2 = "98CCE667333331999999999993333326664CC99B3266CD9B364C9B264D926C9B64DB249B6C9249B6DB6DB6DB692496DB492DA4B692D25A5B4B4B4B4B4A5A5AD296B5AD294A52B5AD4AD6A56A56AD4A952A55AB54AB55AAD56AA554AAB554AAAD5552AAAA5555556AAAAAAAAAAAAAAAAAAAAAAAAAA9555555AAAAB5555AAA9556AA9552AB552A954AB55AB54A952A54A95A952B5295A94AD6B5A94A5AD6B4A52D696B4B4B5A5A5A5B4B4B696D2DA4B692DB492DB692492DB6DB6DB6DB6C924936D924DB24DB24D936C9B26C9B364C9B366CD9B3664CD99332666CCCD9999B33333333333333333333199998CCCE66333998CC673398CE63398C6339CE739CE739";
defparam ram_block1a6.mem_init1 = "CE318E718E718E31C738E39C71C71C71C71C71C70E38F1C78E1C78F1E3C78F1E1C3C7878F0F0F0F0F0F0F078783C3E1F0F83C1F0F83E0F83E07C1F83F07E07E07E07E07E03F81FC07F00FE01FC03FC01FF00FFC01FF801FFC007FF8007FFE0007FFF80003FFFF800000FFFFFFFC0000000000000FFFFFFFFFFFF00000000000001FFFFFFF8000007FFFF80003FFFE0007FFE000FFF8007FF001FF801FF803FF007F803FC03FE03FC03F80FF01FC0FE03F01F80FC0FC0FC0FC0FC1F81F03E0FC1F07E0F83E0F83E1F07C1E0F87C3E1F0F8783C3E1E1F0F0F0F0F8787870F0F0F0E1E1E3C3C7870F1E3C3870E1C3870E3C78E1C78E1C78E3C71E38E1C71C78E38E";
defparam ram_block1a6.mem_init0 = "38E3871C71C718E38E38E38C71C738E39C71CE39C738E71CE31C639C639C631CE318E738C6318E739CE739CE739CE739CE6318CE7398C67398CE7319CC67319CC67319CCE63319CCE673399CCE6633199CCC667331998CCC66633339998CCCC666673333199999CCCCCCCE66666666733333333333333333333333333333333333333333326666666664CCCCCCC999999B33333666664CCCC9999933336666CCCD999B3336666CCC999B332664CCD99B332664CC999332664CD99B33664CC99B32664CD9933666CC99B3266CC9933664CD993366CC99B3664CD9B3264CD9B3264CD9B3264CD9B3664C99B366CC993266CD9B3264C99B366CD993264C99B366CC";

cyclonev_ram_block ram_block1a30(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.clk0_output_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "rom";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "clock0";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 8192;
defparam ram_block1a30.port_a_first_bit_number = 6;
defparam ram_block1a30.port_a_last_address = 16383;
defparam ram_block1a30.port_a_logical_ram_depth = 65536;
defparam ram_block1a30.port_a_logical_ram_width = 24;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init3 = "FFFFFFFFFF00007FFC007FE01FE01FC0FE07C0F83E0F83C1E1E1E1E1C3C78E1C70E38E38C71CE31CE739CE7319CCE6733319999999999333266CC99326CD936C9B6C926DB6DB6DA492DA4B69696D69696B5A5294AD6A56A56AD52AD52AB552AA95552AAAAAB5555555556AAAAAA5554AAA556AA55AA54A952B52B5A94A52D694B4B4B4B4B692DB492DB6DB6DB24936C9B64D9326CD99336664CCCCCCCCCCCCE6673399CC6339CE718C738E31C71C71C38E1C3870F0E1E1F0F0783E0F83F07E07F01FC03FC01FF8007FFE00000FFFFFFFFFFFFFFFC00003FFF000FFC01FF01FE03F03F03E07C1E0F87C3C3C3C3878F1E3871C38E38C71C639C631CE6319CC6733";
defparam ram_block1a30.mem_init2 = "999CCCCCCCCCCCCCC999B3264C99366C93649B64926DB6DB4924B6925A4B4B4B4B4B5A5294A5295A95A952A54AB55AA9552AAD5556AAAAAA955555556AAAAAA95556AAB556AA55AA55AB56A56A52B5AD6B5A52D2D2D2D2DA5B492DB4924924926DB649B24D9366C9933664CC9999993333999998CCE673398C6739CE318E71CE38E38E38E1C78F1E3C387878783C1E0F83E0FC1F80FC07F01FF007FC003FFE0000FFFFFFFFE0003FFFFFFFF80003FFE003FF007F807F01F80FC1F83E0F83C1E0F0F0F0F0E1C3870E38F1C71C738E31C631CE739CC63319CCE667333333333333336664CD9B366CD9364DB26DB249B6DB6DB6924B6D25A4B4969694B4A5AD6B5A";
defparam ram_block1a30.mem_init1 = "D6A56A56A54A956A954AAD55AAAD5556AAAAAA9555555552AAAAAA95556AAB554AAD52A952AD5A95A95A94A5294A5AD2D6969692D25A496D24925B6DB64926DB24D926C99366CD9B32666CCCCD9999998CCCCE6673398CE6319CE738C738C71CE38E38E3C71E3870E1E1C3C3C3E1E0F07C1F07C0F81FC0FE03F807FC01FF8007FFE00003FFFFFFFFFFFFFFFFFFFF80000FFFC007FF007FC03F80FE03F03F07C0F83E1F0F8783C3C7878F0E1C38E1C71C71C71C738E718E739CE7398CE633198CCC666666666666666CCC9993366CD9326C9B64DB24DB6C924924924B6DA4B692DA5A5A5A5A5AD296B5AD6B5A95A95A952A54AB55AAD54AA9554AAA9555552AAA";
defparam ram_block1a30.mem_init0 = "AAAAAAAAAAAAB555556AAAD556AAD54AAD52AD5AB56AD4AD4A56B5AD6B4A52D2D6969692D25A4B6D24B6DB6DB6DB6DB249B649B26D9B26CD9B366CCD99B333326666666733331998CC663398CE739CE739C639C738E38E38E38E3871E3C78F1E1E3C3C3C1E1F0F83C1F03E0FC0FC0FC07F01FE01FF007FF000FFF80003FFFFFE000000000000000FFFFFF80003FFF001FFC00FF007F00FE03F03F03F07E0F83E0F0783C3E1E1E1E3C3878F1E3871C78E38E38E39C718E718E739CE739CC63319CCE663331999999CCCC999999B333666CC993264D9B26C9B24D926DB24936DB6DB6DB4924B6925B4B696D2D2D2D2D696B4A5294A5294AD4A54AD4A952A55AA55";

cyclonev_ram_block ram_block1a103(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a103_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a103.clk0_core_clock_enable = "ena0";
defparam ram_block1a103.clk0_input_clock_enable = "ena0";
defparam ram_block1a103.clk0_output_clock_enable = "ena0";
defparam ram_block1a103.data_interleave_offset_in_bits = 1;
defparam ram_block1a103.data_interleave_width_in_bits = 1;
defparam ram_block1a103.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a103.init_file_layout = "port_a";
defparam ram_block1a103.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a103.operation_mode = "rom";
defparam ram_block1a103.port_a_address_clear = "none";
defparam ram_block1a103.port_a_address_width = 13;
defparam ram_block1a103.port_a_data_out_clear = "none";
defparam ram_block1a103.port_a_data_out_clock = "clock0";
defparam ram_block1a103.port_a_data_width = 1;
defparam ram_block1a103.port_a_first_address = 32768;
defparam ram_block1a103.port_a_first_bit_number = 7;
defparam ram_block1a103.port_a_last_address = 40959;
defparam ram_block1a103.port_a_logical_ram_depth = 65536;
defparam ram_block1a103.port_a_logical_ram_width = 24;
defparam ram_block1a103.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a103.ram_block_type = "auto";
defparam ram_block1a103.mem_init3 = "CCE66331998CCC6666333333199999999999999999933333366664CCD99933266CC99B3264C993264C9B364D9B26C9B26C9364DB26D926D924DB24936DB24924936DB6DB6DB6924924B6DB4925B6925B496D25B496D2DA5B4B4B696969696969694B4B5A5AD296B4A52D6B5AD294AD6B5AD4A52B5295A95A95A95A952B56AD4A952AD5AA54AB54AA55AAD56AA552AB556AAD55AAA5552AAB5552AAAD5554AAAAA555555AAAAAAAA955555555555555555555555555555554AAAAAAAAD555556AAAAB55552AAAD555AAA9554AAB554AA955AAB552A955AAD52A956A956A956AD52A54A952B56AD4AD5A95A95A95AD4AD6A52B5AD4A5294A5294A52D6B4A52D694";
defparam ram_block1a103.mem_init2 = "B5A5AD2D69696B4B4B4B4B4B4969696D2DA5A4B696D25B496D25B692DB4925B6D2492DB6DA4924924924924924924DB6DB24926DB64936C926D926D926C93649B26C9B64D9326C9B264D9326CD9B264C993366CD9933664CD99B32666CCD999B333666664CCCCCD999999999999999999999999998CCCCCC666673333999CCCE66733198CCE673398CC673398CE63398C67318CE7398C6318C6318C6318C631CE718C738C639C638C738E71CE39C718E38C71C718E38E38E38E38E38E38E3871C71C38E3C71C38F1C78E1C78F1C3870E1C3870E1C3C78F0E1E1C3C387878F0F0F0F0F0F0F0F0F0F0F8787C3C3E1E0F0787C3E0F0783E1F07C3E0F83E0F83E0F8";
defparam ram_block1a103.mem_init1 = "3E0F81F07E0F81F03F07E07C0FC0FC0FC0FC0FC07E07F03F81FC07F01FC07F01FC03F807F00FF00FF00FF007F803FE00FF803FF007FE007FF003FF800FFE001FFE001FFF0007FFC000FFFE0003FFFE0000FFFFC00007FFFFC000007FFFFFE00000007FFFFFFFFC0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000FFFFFFFFFC00000007FFFFFF000000FFFFFE00001FFFFC00007FFFC0003FFFC0003FFF0001FFF0003FFE000FFF000FFF000FFE003FF800FFE007FF003FF003FE007FC00FF803FE00FF803FC01FE00FF00FF007F80FF00FF00FE01FC03F807F01FC07F80FE03F80FC07F01F80FE07F03F81FC0FC07E07F03F0";
defparam ram_block1a103.mem_init0 = "3F03F01F81F83F03F03F03E07E07C0FC1F81F03E07C0F81F03E07C1F83E07C1F03E0F83E07C1F07C1F07C1F07C1F07C1F07C1F0F83E0F87C1F0F83E1F0783E1F0783E1F0F83C1E0F0783C1E0F0783C1E1F0F8783C1E1F0F0787C3C3E1E0F0F078787C3C3C1E1E1F0F0F0F0787878787C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C387878787878F0F0F0E1E1E1E3C3C3C787878F0F0E1E1C3C3C7878F0F1E1E3C3C7878F0F1E1C3C7878F0E1E3C387870F1E1C3C78F0E1E3C3878F0E1C3C7870E1E3C7870E1E3C3870E1E3C7870E1E3C78F0E1C3878F1E3C3870E1C3C78F1E3C3870E1C3878F1E3C78F0E1C3870E1C3C78F1E3C78F1E1C3870E1C3870E";

cyclonev_ram_block ram_block1a127(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a127_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a127.clk0_core_clock_enable = "ena0";
defparam ram_block1a127.clk0_input_clock_enable = "ena0";
defparam ram_block1a127.clk0_output_clock_enable = "ena0";
defparam ram_block1a127.data_interleave_offset_in_bits = 1;
defparam ram_block1a127.data_interleave_width_in_bits = 1;
defparam ram_block1a127.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a127.init_file_layout = "port_a";
defparam ram_block1a127.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a127.operation_mode = "rom";
defparam ram_block1a127.port_a_address_clear = "none";
defparam ram_block1a127.port_a_address_width = 13;
defparam ram_block1a127.port_a_data_out_clear = "none";
defparam ram_block1a127.port_a_data_out_clock = "clock0";
defparam ram_block1a127.port_a_data_width = 1;
defparam ram_block1a127.port_a_first_address = 40960;
defparam ram_block1a127.port_a_first_bit_number = 7;
defparam ram_block1a127.port_a_last_address = 49151;
defparam ram_block1a127.port_a_logical_ram_depth = 65536;
defparam ram_block1a127.port_a_logical_ram_width = 24;
defparam ram_block1a127.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a127.ram_block_type = "auto";
defparam ram_block1a127.mem_init3 = "000000000000007FFFFF80001FFFE000FFF800FFC00FFC01FE01FE01FC07F01F81FC0FC0F81F03E0F83E0F83E1F0F87C3C3E1E1E1E1E1C3C3870F1E3C70E1C70E38F1C71C71C71C718E38C718E718E718C639CE7318C67398CE63319CCC6633319998CCCCCC6666666664CCCCCD9999332664CC993366CD9B264D9326C9B64D926D926D924DB6D92492492492492DB6D2496DA4B692DA5B4B4969696969696B4B5A52D6B4A5294A5295AD4A56A56A56AD5A952A55AA54AA55AAD54AAD55AAB555AAA95556AAAAD555555AAAAAAAAAAAAAAAAAAAAAAAAA9555555AAAAB5554AAAD556AA955AAB55AAD56A956A952A54A952B52A56A52B5294AD6B5AD6B4A52D69";
defparam ram_block1a127.mem_init2 = "4B4A5A5A5A5A5A5A5B4B696D25B492DB492DB6D24924924924926DB64926D926D926C9364D9366C9B364C993266CC99B336664CCCD9999999333333319999998CCCE66733199CC663398CE6319CE739CE739CE31CE31CE39C738E38C71C71C71E38E3871C38F1E3870F1E3C38787878F0F878787C3E1F0F87C1F07C1F07E0FC1F81F81F80FC07F01FC07F807FC03FE007FE003FF8003FFF0000FFFFE000001FFFFFFFFFFFFF801FFFFFFFFFFFFFC000003FFFF80007FFE000FFE003FF003FE00FF00FF01FE03F81FC0FE07E07C0FC1F83E0F83E0F87C1E0F0787C3C3C3C3C3C3C3878F0E1C3870E1C78E3C71C38E38E38E38E38C71C638C738E738C739CE739C";
defparam ram_block1a127.mem_init1 = "E7398C67398CE673198CCE6633319998CCCCCCC66666666CCCCCCC9999B332664CC99B3264C99326CD9326C9B26C93649B24DB249B6D924936DB6DB6DB6DB492496DA496DA4B692DA4B4B69696D2D2D2D69694B4A5AD294B5AD6B5AD6A5295A94AD4AD4A95AB52A55AB56A956AB54AA556AA556AA9556AAB5552AAA955556AAAAAB555555555555555555555555555554AAAAAAD55552AAA9555AAA9556AAD55AA954AA552AD56AD52A55AB52A54AD4AD4AD4AD6A52B5AD6B5AD6B5A5296B4A5A5AD2D2D2D2D2D2D25A5B4B692DA4B6D25B6D2496DB6DA4924924936DB6D9249B6C936C936C9B64D9364D9364C9B364C993366CC99B32664CCD9999333336666";
defparam ram_block1a127.mem_init0 = "6666666666667333331999CCCE6633399CCE63398CE6339CC6318C6318C639CE318E71CE31C638E31C71C71C71C71C71C78E3871E3871E3C78F1E3C3878F0F0F1E1E1E1F0F0F0787C3E1F0783E0F83E0F83E07C0F81F81F81F81FC0FE03F80FE01FC03FE01FF007FC00FFE003FFC003FFF0001FFFF00000FFFFFF80000000001FFFFFFFFFFFFFFF00000000003FFFFFE00001FFFF8000FFF8003FFC007FF003FF007FC03FE01FE03FC07F01FC07E07F03F03F03E07E0F81F07C1F07C1F0783E1F0F87C3C1E1E1E1F0F1E1E1E1C3C3878F1E1C3871E3C70E3C71E38E3C71C71C71C71C71C638E39C738E71CE31CE318E738C6318C6318CE7318CE7319CC663399";

cyclonev_ram_block ram_block1a151(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a151_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a151.clk0_core_clock_enable = "ena0";
defparam ram_block1a151.clk0_input_clock_enable = "ena0";
defparam ram_block1a151.clk0_output_clock_enable = "ena0";
defparam ram_block1a151.data_interleave_offset_in_bits = 1;
defparam ram_block1a151.data_interleave_width_in_bits = 1;
defparam ram_block1a151.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a151.init_file_layout = "port_a";
defparam ram_block1a151.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a151.operation_mode = "rom";
defparam ram_block1a151.port_a_address_clear = "none";
defparam ram_block1a151.port_a_address_width = 13;
defparam ram_block1a151.port_a_data_out_clear = "none";
defparam ram_block1a151.port_a_data_out_clock = "clock0";
defparam ram_block1a151.port_a_data_width = 1;
defparam ram_block1a151.port_a_first_address = 49152;
defparam ram_block1a151.port_a_first_bit_number = 7;
defparam ram_block1a151.port_a_last_address = 57343;
defparam ram_block1a151.port_a_logical_ram_depth = 65536;
defparam ram_block1a151.port_a_logical_ram_width = 24;
defparam ram_block1a151.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a151.ram_block_type = "auto";
defparam ram_block1a151.mem_init3 = "3398CC67319CE6319CE6318C6318C639CE318E718E71CE39C738E38C71C71C71C71C71C78E38F1C78E1C78F1C3870F1E3C387870F0F0F1E1F0F0F0F0787C3E1F0F83C1F07C1F07C1F03E0FC0F81F81F81FC0FC07F01FC07F80FF00FF807FC01FF801FFC007FF8003FFE0003FFFF00000FFFFFF80000000001FFFFFFFFFFFFFFF00000000003FFFFFE00001FFFF0001FFF8007FF800FFE007FC01FF00FF807F00FE03F80FE07F03F03F03F03E07C0F83E0F83E0F83C1F0F87C3C1E1E1F0F0F0F1E1E1E3C3878F1E3C78F1C38F1C38E3C71C71C71C71C71C718E38C718E71CE318E738C6318C6318C67398CE63398CE6733998CCE667333199999CCCCCCCCCCCCC";
defparam ram_block1a151.mem_init2 = "CCCD9999933336664CC99B3266CD993264D9B264D9364D9364DB26D926D926DB24936DB6D924924924B6DB6D2496DB496DA4B692DA5B4B496969696969696B4B4A5AD294B5AD6B5AD6B5A94AD6A56A56A56A54A95AB54A956AD56A954AA552AB556AAD552AAB5552AAA955556AAAAAA555555555555555555555555555555AAAAAAD55552AAA9555AAAD552AAD54AAD54AA55AAD52AD5AB54A95AB52A56A56A52B5294AD6B5AD6B5A5296B4A5A52D2D6969696D2D2DA5A4B692DA4B6D24B6D24925B6DB6DB6DB6D924936DB249B649B24D926C9B26C99366C993264C99B32664CC999B33326666666CCCCCCCC666666633331998CCE663319CCE6339CC6339CE";
defparam ram_block1a151.mem_init1 = "739CE739C639CE39C638C71C638E38E38E38E3871C78E3C70E1C3870E1E3C387878787878787C3C1E0F07C3E0F83E0F83F07E07C0FC0FE07F03F80FF01FE01FE00FF801FF800FFE000FFFC0003FFFF8000007FFFFFFFFFFFFF003FFFFFFFFFFFFF000000FFFFE0001FFF8003FF800FFC00FF807FC03FC07F01FC07E03F03F03F07E0FC1F07C1F07C3E1F0F87C3C3C3E1E3C3C3C3878F1E1C38F1E3871C38E38F1C71C71C638E39C738E718E718E739CE739CE7318CE63398CC6733199CCCE666333333319999999333333366664CCD99B3266CC993264D9B26CD9364D926C936C936C924DB6C92492492492496DB6925B6925B496D2DA5B4B4B4B4B4B4B4A5A5";
defparam ram_block1a151.mem_init0 = "2D694A5AD6B5AD6A5295A94AD4A95A952A54A952AD52AD56AB55AAB552AAD556AAA5555AAAAB5555552AAAAAAAAAAAAAAAAAAAAAAAAB5555556AAAAD5552AAB555AAB556AA556AB54AA54AB54A952B56AD4AD4AD4A56B5294A5294A5AD694B5A5AD2D2D2D2D2D25A5B4B692DA4B6D2496DB6924924924924936DB64936C936C9364DB26C99364C9B366CD9932664CC99933336666664CCCCCCCCC66666633331998CC6673198CE6339CC6319CE738C631CE31CE31C638E31C71C71C71C71E38E1C70E1C78F1E1C387870F0F0F0F0F8787C3E1F0F83E0F83E0F81F03E07E07F03F01FC07F00FF00FF007FE007FE003FFE000FFFF00003FFFFFC00000000000000";

cyclonev_ram_block ram_block1a175(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a175_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a175.clk0_core_clock_enable = "ena0";
defparam ram_block1a175.clk0_input_clock_enable = "ena0";
defparam ram_block1a175.clk0_output_clock_enable = "ena0";
defparam ram_block1a175.data_interleave_offset_in_bits = 1;
defparam ram_block1a175.data_interleave_width_in_bits = 1;
defparam ram_block1a175.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a175.init_file_layout = "port_a";
defparam ram_block1a175.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a175.operation_mode = "rom";
defparam ram_block1a175.port_a_address_clear = "none";
defparam ram_block1a175.port_a_address_width = 13;
defparam ram_block1a175.port_a_data_out_clear = "none";
defparam ram_block1a175.port_a_data_out_clock = "clock0";
defparam ram_block1a175.port_a_data_width = 1;
defparam ram_block1a175.port_a_first_address = 57344;
defparam ram_block1a175.port_a_first_bit_number = 7;
defparam ram_block1a175.port_a_last_address = 65535;
defparam ram_block1a175.port_a_logical_ram_depth = 65536;
defparam ram_block1a175.port_a_logical_ram_width = 24;
defparam ram_block1a175.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a175.ram_block_type = "auto";
defparam ram_block1a175.mem_init3 = "E1C3870E1C3870F1E3C78F1E3C7870E1C3870E1E3C78F1E3C3870E1C3878F1E3C7870E1C3878F1E3C3870E1E3C78F0E1C3C78F0E1C3878F0E1C3C78F0E1C3C7870E1E3C3878F0E1E3C7870F1E1C3C3878F0E1E3C3C7870F1E1E3C3C7878F0F1E1E3C3C787870F0E1E1E3C3C3C787878F0F0F0E1E1E1E3C3C3C3C3C3878787878787878787878787878787878787878787C3C3C3C3C1E1E1E1F0F0F078787C3C3C1E1E0F0F8787C3C1E1F0F0783C3E1F0F0783C1E0F0783C1E0F0783E1F0F83C1F0F83C1F0F83E1F07C3E0F83E1F07C1F07C1F07C1F07C1F07C1F07C0F83E0F81F07C0F83F07C0F81F03E07C0F81F03F07E07C0FC0F81F81F81F83F03F01F81F8";
defparam ram_block1a175.mem_init2 = "1F81FC0FC07E07F03F81FC0FE03F01FC07E03F80FE03FC07F01FC03F807F00FE01FE01FE03FC01FE01FE00FF007F803FE00FF803FE007FC00FF801FF801FFC00FFE003FF800FFE001FFE001FFE000FFF8001FFF0001FFF80007FFF80007FFFC00007FFFF00000FFFFFE000001FFFFFFC00000007FFFFFFFFE00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000007FFFFFFFFC0000000FFFFFFC000007FFFFC00007FFFE0000FFFF8000FFFE0007FFC001FFF000FFF000FFE003FF801FFC00FFC01FF803FE00FF803FC01FE01FE01FE01FC03F807F01FC07F01FC07F03F81FC0FC07E07E07E07E07E07C0FC1F81F03E0FC1F03E0F8";
defparam ram_block1a175.mem_init1 = "3E0F83E0F83E0F87C1F0F83C1E0F87C3C1E0F0F8787C3C3E1E1E1E1E1E1E1E1E1E1E3C3C387870F0E1E3C7870E1C3870E1C3871E3C70E3C71E3871C78E3871C71C38E38E38E38E38E38E38E31C71C638E31C738E71CE39C638C738C639C631CE718C6318C6318C6318C6339CE6319CC63398CE63399CC663399CCE6633199CCCE6673339999CCCCC6666663333333333333333333333333336666664CCCCD999B333666CCC99B33664CD993366CD993264C9B366C99364C9B26C99364DB26C9B24D926C936C936C926D924DB6C9249B6DB64924924924924924924B6DB692496DB4925B692DB496D25B496D2DA4B4B696D2D2D25A5A5A5A5A5AD2D2D696B4B5A";
defparam ram_block1a175.mem_init0 = "52D694A5AD694A5294A5294A56B5A94AD6A56B52B52B52B56A56AD5A952A54A956AD52AD52AD52A956AB552A955AAB552AA555AAA5552AAB5556AAA95555AAAAAD555556AAAAAAAA555555555555555555555555555555552AAAAAAAB555554AAAAA55556AAA9555AAA9554AAB556AAD55AA954AAD56AB54AA55AA54AB56A952A56AD5A952B52B52B52B5295A94A56B5AD6A5296B5AD694A5AD296B4B5A5A52D2D2D2D2D2D2DA5A5B4B696D25B496D25B492DB4925B6DA492492DB6DB6DB6D9249249B6D9249B64936C936C9B64D926C9B26C9B364D9B264C993264C99B3266CC9993336664CCCD9999993333333333333333331999998CCCC666333198CCE67";

cyclonev_ram_block ram_block1a55(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a55_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a55.clk0_core_clock_enable = "ena0";
defparam ram_block1a55.clk0_input_clock_enable = "ena0";
defparam ram_block1a55.clk0_output_clock_enable = "ena0";
defparam ram_block1a55.data_interleave_offset_in_bits = 1;
defparam ram_block1a55.data_interleave_width_in_bits = 1;
defparam ram_block1a55.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a55.init_file_layout = "port_a";
defparam ram_block1a55.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a55.operation_mode = "rom";
defparam ram_block1a55.port_a_address_clear = "none";
defparam ram_block1a55.port_a_address_width = 13;
defparam ram_block1a55.port_a_data_out_clear = "none";
defparam ram_block1a55.port_a_data_out_clock = "clock0";
defparam ram_block1a55.port_a_data_width = 1;
defparam ram_block1a55.port_a_first_address = 16384;
defparam ram_block1a55.port_a_first_bit_number = 7;
defparam ram_block1a55.port_a_last_address = 24575;
defparam ram_block1a55.port_a_logical_ram_depth = 65536;
defparam ram_block1a55.port_a_logical_ram_width = 24;
defparam ram_block1a55.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a55.ram_block_type = "auto";
defparam ram_block1a55.mem_init3 = "CC673398CE6319CC6319CE739CE739C631CE718E718E31C638C71C638E38E38E38E38E3871C70E3871E3870E3C78F1E1C3C7878F0F0F1E1E0F0F0F0F8783C1E0F0783E0F83E0F83E0FC1F03F07E07E07E03F03F80FE03F807F00FF007F803FE007FE003FF8007FF8001FFFC0001FFFFF0000007FFFFFFFFFE000000000000000FFFFFFFFFFC000001FFFFE0000FFFE0007FF8007FF001FF803FE00FF807F80FF01FC07F01FC0FC0FC0FC0FC1F83F07C1F07C1F07C3E0F0783C3E1E1E0F0F0F0F1E1E1C3C7870E1C3870E3C70E3C71C38E38E38E38E38E38E71C738E71CE31CE718E739CE739CE7398C67319CC673198CC667331998CCCE666663333333333333";
defparam ram_block1a55.mem_init2 = "3332666664CCC999B33664CD993366CD9B264D9B26C9B26C9B24D926D926D924DB6C924936DB6DB6DB492492DB6924B6D25B496D25A4B4B696969696969696B4B5A52D6B4A5294A5294A56B5295A95A95A95AB52A54AB56A952AD56AB55AAD54AA9552AAD554AAAD5556AAAA9555554AAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5555556AAAAD5556AAA5552AA9552AB552AB55AA552AD52A55AB56A54AD5A95A95AD4AD6B5294A5294A5AD694B5A5AD2D296969692D2D25A5B496D25B496DA492DB6DA4924924924924DB6D924DB649B64DB26D9364D9366C99366CD9B3664CD993336664CCC9999999B333333331999999CCCCE66733199CCE63319CC6339CC631";
defparam ram_block1a55.mem_init1 = "8C6318C639CE31CE39C738E39C71C71C71C71C78E3871C38F1E3C78F1E3C3C787878787878783C3E1F0F87C1F07C1F07C0F81F83F03F01F81FC07F01FE01FE01FF007FE007FF001FFF0003FFFC00007FFFFF80000000000007FFF0000000000000FFFFFF80001FFFE0007FFC007FF003FF007FC03FC03F80FE03F80FC0FC0FC0F81F03E0F83E0F83C1E0F0783C3C3C1E1E3C3C3C7870E1E3C70E1C78E3C71C70E38E38E39C71C638C718E718E718C6318C6318CE7319CC673398CCE663331999CCCCCCCE66666664CCCCCC9999B332664CD993366CD9B264D9B26C9B26D936C936C936D924936DB6DB6DB6DB692496DB496DA4B692D25A4B4B4B4B4B4B4B5A5A";
defparam ram_block1a55.mem_init0 = "D296B5A5294A5295AD6A56B52B52A56AD5AB56AD52AD52A954AA556AAD552AAD555AAAA55554AAAAAAD5555555555555555555555555AAAAAA955552AAAD554AAA554AA955AA954AB55AA54AB56AD5A952B52B52B5A94AD6B5AD6B5AD296B4A5A52D2D2D2D2D2D25A4B496D25B492DB6924B6DB6DB6DB6DB6C9249B6C936C936C9B24D9366C9B364C993266CD99B32666CCCD999999B3333333339999998CCCE66733998CE67319CC6339CE6318C739CE31CE31CE39C718E38E38E38E38E1C71E38F1E3870E1E3C7878F0F0F0F0F0F8783C1E0F07C1F07C1F07E0FC1F81F81FC0FE03F80FF00FF00FF801FF801FFC001FFF0000FFFFC000003FFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a79(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a79_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a79.clk0_core_clock_enable = "ena0";
defparam ram_block1a79.clk0_input_clock_enable = "ena0";
defparam ram_block1a79.clk0_output_clock_enable = "ena0";
defparam ram_block1a79.data_interleave_offset_in_bits = 1;
defparam ram_block1a79.data_interleave_width_in_bits = 1;
defparam ram_block1a79.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a79.init_file_layout = "port_a";
defparam ram_block1a79.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a79.operation_mode = "rom";
defparam ram_block1a79.port_a_address_clear = "none";
defparam ram_block1a79.port_a_address_width = 13;
defparam ram_block1a79.port_a_data_out_clear = "none";
defparam ram_block1a79.port_a_data_out_clock = "clock0";
defparam ram_block1a79.port_a_data_width = 1;
defparam ram_block1a79.port_a_first_address = 24576;
defparam ram_block1a79.port_a_first_bit_number = 7;
defparam ram_block1a79.port_a_last_address = 32767;
defparam ram_block1a79.port_a_logical_ram_depth = 65536;
defparam ram_block1a79.port_a_logical_ram_width = 24;
defparam ram_block1a79.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a79.ram_block_type = "auto";
defparam ram_block1a79.mem_init3 = "1E3C78F1E3C78F0E1C3870E1C3878F1E3C78F1E1C3870E1C3C78F1E3C7870E1C3878F1E3C7870E1C3C78F1E1C3870F1E3C3870E1E3C7870E1E3C3870F1E3C3878F1E1C3C7870F1E3C3878F0E1E3C387870F1E1C3C7878F0E1E1C3C387870F0E1E1C3C387870F0F1E1E1C3C3C38787870F0F0E1E1E1E1C3C3C3C3C387878787878787878787878787878787878787878783C3C3C3C3E1E1E1E0F0F0F078783C3C3E1E1F0F078783C3E1E0F0F87C3C1E0F0F87C3E1F0F87C3E1F0F87C1E0F07C3E0F07C3E0F07C1E0F83C1F07C1E0F83E0F83E0F83E0F83E0F83E0F83E07C1F07E0F83F07C0F83F07E0FC1F83F07E0FC0F81F83F03E07E07E07E0FC0FC0FC07E07";
defparam ram_block1a79.mem_init2 = "E07E03F03F01F80FC07E03F01FC0FE03F81FC07F01FC07F80FE03FC07F80FF01FE01FE03FC03FE01FE01FF00FF807FC01FF007FC01FF003FF007FE007FE003FF001FF800FFF001FFE001FFE001FFF0007FFE000FFFE0007FFF80007FFF80003FFFF80000FFFFF000003FFFFFE0000003FFFFFFF8000000003FFFFFFFFFFFFF0000000000000000000000000000000000000007FFFFFFFFFFFFC000000003FFFFFFF0000003FFFFF800003FFFF80001FFFF80007FFF0001FFF8003FFF000FFF000FFF001FFC007FF003FF003FE007FC01FF007FC03FE01FE01FE01FE03FC07F80FE03F80FE03F80FC07E03F01F81F81F81F81F81F83F03E07E0FC1F03E0FC1F07";
defparam ram_block1a79.mem_init1 = "C1F07C1F07C1F07C3E0F07C3E1F0783C3E1F0F0787C3C3C1E1E1E1E1E1E1E1E1E1E1C3C3C7878F0F1E1C3878F1E3C78F1E3C78E1C38F1C38E1C78E3871C78E38E1C71C71C71C71C71C71C71CE38E39C71CE38C718E31C639C738C739C639CE318E739CE738C6339CE739CC6319CE6339CC67319CC663399CC6633199CCE66333199CCCC666633333999999CCCCCCCCCCCCCCCCCCCCCCCCCCC9999999333326664CCC999333666CC99B3266CC993266CD9B364C99366C9B364D9326C9B24D9364DB26D936C936C936D926DB24936DB249249B6DB6DB6DB6DB6DB6DB492492DB6924B6DA496D24B692DA4B692D25B4B69692D2D2DA5A5A5A5A5A52D2D29694B4A5";
defparam ram_block1a79.mem_init0 = "AD296B5A5296B5AD6B5AD6B5A94A56B5295AD4AD4AD4AD4AD5A952B56AD5AB56A952AD52AD52AD56A954AAD56AA556AAD55AAA555AAAD554AAA95556AAAA555552AAAAA955555554AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAD55555554AAAAAA55555AAAA95556AAA5556AAB554AA9552AA556AB552A954AB55AA55AB54A956AD5AB52A56AD4AD4AD4AD4AD6A56B5A94A52B5AD694A5296B5A52D694B4A5A5AD2D2D2D2D2D2D25A5A4B49692DA4B492DA4B6D24B6DA4925B6DB6924924924924DB6DB64926DB649B6C936C93649B26D9364D9364C9B264D9B366CD9B3664CD9933666CCC999B3332666666CCCCCCCCCCCCCCCCCCE6666673333999CCCE6633198";

cyclonev_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 8191;
defparam ram_block1a7.port_a_logical_ram_depth = 65536;
defparam ram_block1a7.port_a_logical_ram_width = 24;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init3 = "33198CCE6673339999CCCCCCE666666666666666666CCCCCC9999B332666CCD9933664CD9B366CD9B364C9B264D9364D936C9B24D926D926DB24DB6C924DB6DB6492492492492DB6DB4924B6DA496DA4B6925A4B692D25A4B4B496969696969696B4B4A5A52D694B5AD294A52D6B5A94A52B5AD4AD6A56A56A56A56AD4A95AB56AD52A55AB54AB55AA552A955AAD54AA9552AA555AAAD554AAAD5552AAAB55554AAAAAA555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA555555552AAAAA955554AAAAD5552AAA5556AAB554AAB556AAD54AAD56AA552AD56A956A956A952AD5AB56AD5A952B56A56A56A56A56B5295AD4A52B5AD6B5AD6B5AD294B5AD296B";
defparam ram_block1a7.mem_init2 = "4A5A52D2969694B4B4B4B4B4B6969692D2DA5B49692DA4B692DA496D24B6DA492DB6924925B6DB6DB6DB6DB6DB6DB249249B6D9249B6C936D926D926D936C9B64D93649B26C99364D9B26CD93264D9B366CC993266CC99B3266CCD9993326664CCC99999333333266666666666666666666666666733333399998CCCC6667331998CCE6733198CC673398CC67319CC67398CE7318C6739CE7398C639CE739CE318E738C739C639C738C718E31C638E71C738E38E71C71C71C71C71C71C71C70E38E3C71C38E3C70E3871E3870E3C78F1E3C78F1E3C3870F1E1E3C3C787870F0F0F0F0F0F0F0F0F0F078787C3C1E1F0F8783C1F0F87C1E0F87C1F07C1F07C1F07";
defparam ram_block1a7.mem_init1 = "C1F07E0F81F07E0FC0F81F83F03F03F03F03F03F01F80FC07E03F80FE03F80FE03FC07F80FF00FF00FF00FF807FC01FF007FC00FF801FF801FFC007FF001FFE001FFE001FFF8003FFF0001FFFC0003FFFF00003FFFF800003FFFFF8000001FFFFFFF8000000007FFFFFFFFFFFFC000000000000000000000000000000000000001FFFFFFFFFFFFF8000000003FFFFFFF8000000FFFFFF800001FFFFE00003FFFF80003FFFC0003FFFC000FFFE000FFFC001FFF000FFF000FFF001FFE003FF001FF800FFC00FFC01FF801FF007FC01FF007FC03FE01FF00FF00FF807F80FF00FF01FE03FC07F80FE03FC07F01FC07F03F80FE07F01F80FC07E03F01F81F80FC0F";
defparam ram_block1a7.mem_init0 = "C0FC07E07E07E0FC0FC0FC0F81F83F03E07E0FC1F83F07E0FC1F83E07C1F83E0FC1F07C0F83E0F83E0F83E0F83E0F83E0F83E0F07C1F0783E0F07C1E0F87C1E0F87C1E0F07C3E1F0F87C3E1F0F87C3E1E0F0787C3E1E0F0F8783C3C1E1F0F0F878783C3C1E1E1E0F0F0F0F8787878783C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C3C387878787870F0F0F0E1E1E1C3C3C38787870F0F1E1E1C3C387870F0E1E1C3C387870F0E1E3C3C7870F1E1C3C3878F0E1E3C3878F1E1C3C7870F1E3C3878F1E1C3878F0E1C3C78F0E1C3878F1E1C3870F1E3C7870E1C3C78F1E3C3870E1C3C78F1E3C7870E1C3870F1E3C78F1E3C3870E1C3870E1E3C78F1E3C78F0";

cyclonev_ram_block ram_block1a31(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.clk0_output_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "rom";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "clock0";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 8192;
defparam ram_block1a31.port_a_first_bit_number = 7;
defparam ram_block1a31.port_a_last_address = 16383;
defparam ram_block1a31.port_a_logical_ram_depth = 65536;
defparam ram_block1a31.port_a_logical_ram_width = 24;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init3 = "FFFFFFFFFFFFFF8000007FFFE0001FFF0007FF003FF003FE01FE01FE03F80FE07F03F03F07E0FC1F07C1F07C1E0F0783C3E1E1E1E1E1E3C3C78F0E1C38F1E38F1C70E38E38E38E38E31C738E718E718E739C6318CE7398C67319CCE633399CCCE6663333333999999999B3333336666CCC99B3366CC993264D9B26CD93649B26D926D926DB24926DB6DB6DB6DB6DA492DB6925B496D25A4B496969696969694B4A5AD296B5AD6B5AD6A52B5A95A95A952B56AD5AA54AB55AA552AB552AA554AAA5556AAA955552AAAAAB55555555555555555555555556AAAAAA55554AAAB5556AA9556AAD54AA552A956A956AD5AB56AD4A95A95AD4AD6B5294A5294B5AD296";
defparam ram_block1a31.mem_init2 = "B4B5A5A5A5A5A5A5A4B49692DA4B6D25B6D2492DB6DB6DB6DB6D924936D926D926D936C9B26C9B364C9B366CD9933664CC999B33326666664CCCCCCCE66666673331998CCE663399CC67319CE6318C6318C631CE31CE31C638C71C738E38E38E1C71C78E3C70E1C78F0E1C3C787878F0F07878783C1E0F0783E0F83E0F81F03E07E07E07E03F80FE03F807F807FC01FF801FFC007FFC000FFFF00003FFFFFE0000000000001FFFC0000000000003FFFFFC00007FFF8001FFF001FFC00FFC01FF00FF00FF01FC07F03F01F81F83F03E07C1F07C1F07C3E1F0F8783C3C3C3C3C3C3C7878F1E3C78F1E3871C38E3C71C71C71C71C738E39C738E718E738C6318C63";
defparam ram_block1a31.mem_init1 = "18C67398C673198CE6733199CCCE6667333333199999999B33333326664CCD99933664CD9B366CD9326CD9364D936C9B64DB24DB64936DB64924924924924B6DB6924B6D25B496D25B4B4969692D2D2D29696B4B5A52D6B4A5294A5295AD6A56B52B52B56A54AD5AB54A956A954AB55AA955AA9552AA9554AAAD5556AAAAD555554AAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5555552AAAAD5556AAA5556AA9552AA556AB55AAD56A952AD5AA54A95AB52B52B52B5295AD4A5294A5294A5AD694B5A5AD2D2D2D2D2D2D2DA5A4B496D25B496DA492DB6924925B6DB6DB6D924926DB64936C936C93649B26C9B26C9B364C9B366CD9933664CD99B3326664CCCCC9999";
defparam ram_block1a31.mem_init0 = "9999999999998CCCCCE666333199CCC663319CC67319CC6339CE739CE739CE31CE718E71CE39C71CE38E38E38E38E38E3871C78E1C78E1C3870E1C3C7870F0F1E1E1E1E0F0F0F8783C1E0F87C1F07C1F07C1F83F07E07E07E07E07F01FC07F01FE03FC03FE00FF803FF001FFC003FFC000FFFE0000FFFFF0000007FFFFFFFFFE000000000000000FFFFFFFFFFC000001FFFFF00007FFF0003FFC003FF800FFC00FF803FC01FE01FC03F80FE03F81F80FC0FC0FC1F81F07E0F83E0F83E0F83C1E0F0783C3E1E1E1E0F0F1E1E1E3C3C7870F1E3C78E1C38F1C38E1C71C38E38E38E38E38E38C71C638C718E31CE31CE718C739CE739CE7318C67318CE63399CC66";

cyclonev_ram_block ram_block1a104(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a104_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a104.clk0_core_clock_enable = "ena0";
defparam ram_block1a104.clk0_input_clock_enable = "ena0";
defparam ram_block1a104.clk0_output_clock_enable = "ena0";
defparam ram_block1a104.data_interleave_offset_in_bits = 1;
defparam ram_block1a104.data_interleave_width_in_bits = 1;
defparam ram_block1a104.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a104.init_file_layout = "port_a";
defparam ram_block1a104.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a104.operation_mode = "rom";
defparam ram_block1a104.port_a_address_clear = "none";
defparam ram_block1a104.port_a_address_width = 13;
defparam ram_block1a104.port_a_data_out_clear = "none";
defparam ram_block1a104.port_a_data_out_clock = "clock0";
defparam ram_block1a104.port_a_data_width = 1;
defparam ram_block1a104.port_a_first_address = 32768;
defparam ram_block1a104.port_a_first_bit_number = 8;
defparam ram_block1a104.port_a_last_address = 40959;
defparam ram_block1a104.port_a_logical_ram_depth = 65536;
defparam ram_block1a104.port_a_logical_ram_width = 24;
defparam ram_block1a104.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a104.ram_block_type = "auto";
defparam ram_block1a104.mem_init3 = "C3E1E0F0787C3C1E1E0F0F0F0787878787878787878F0F0F0E1E1C3C3878F0E1E3C7870E1C3870E1C3870E3C78E1C78E1C70E3C71E38E1C71C38E38F1C71C71C70E38E38E38E71C71C71C738E38E71C738E31C738E31C638C738E718E718E718E738C739C6318E739CE318C6318C6318C6339CE7318C67398C67398CE7319CC67319CC663398CC663399CCE6633198CCE66333999CCCE6673331999CCCCC66666333333999999998CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCD99999999B33333266666CCCC9999B3336664CCD999332664CC99933664CC99B3664CD9B3264CD9B366CD9B366CD9B264C9B364C9B364D9B26C99364D9364D9364D9364D926C9B24D";
defparam ram_block1a104.mem_init2 = "936C9B64DB24D926D926D926DB24DB249B6C926DB24936DB24936DB64924936DB6DB6492492492492492492492492492496DB6DB6D24925B6DB4924B6DA492DB6925B6D24B6925B692DB496DA4B692DA4B692DA4B496D2DA4B49692D25A4B4B69692D2D2DA5A5A4B4B4B4B4B4B4B4B4B4B4B4B4B4A5A5A5AD2D2D69694B4A5A52D296B4A5A52D694A5AD296B5A5296B5AD294A5AD6B5AD6B5AD6B5AD6B5AD6B5AD4A5295AD6B5295AD6A52B5A94AD4A56A52B52B5A95A95A95A95A95A95A952B52B56A56AD4A95AB52A54AD5AB56AD5AB56AD5AB56AD5AA54AB56A952AD5AA55AA55AA55AA55AA55AAD52A956AB55AAD52A955AAD56AB552A955AA955AA955AA";
defparam ram_block1a104.mem_init1 = "955AAB552AA554AA9552AAD55AAA555AAA555AAAD552AA9554AAAD554AAAD554AAA95552AAA5555AAAA55552AAA95555AAAA955552AAAAD55556AAAAA555554AAAAAB5555552AAAAAA55555556AAAAAAAA5555555552AAAAAAAAAAD55555555555552AAAAAAAAAAAAAAAAAAAAA9555555555555555555555555555555555555556AAAAAAAAAAAAAAAAAAAAAA955555555555555AAAAAAAAAAAB5555555556AAAAAAAA955555556AAAAAAA5555555AAAAAAB555555AAAAAA555554AAAAAD55554AAAAA55555AAAAB55556AAAAD5554AAAAD5556AAAB5555AAAA55552AAA5555AAAB5556AAAD555AAA95552AAB5552AA9555AAAD554AAA5552AA9556AAB555AAA5";
defparam ram_block1a104.mem_init0 = "55AAA5552AAD55AAA555AAB554AA9556AAD55AAB556AAD55AAB556AAD54AA955AAB552AB556AA556AA556AA556AA556AA556AA552AB552A955AAD54AA552AB55AAD54AA552A954AA552A954AA552A954AA552AD56AB55AA552A956AB54AA55AAD52A956A954AB55AA55AA552AD52AD56A956A956A956A956A956A956A956A956A956A956AD52AD52AD52A55AA54AB54AB56A956AD52AD5AA54AB56A956AD52A55AB54A956AD52A55AB56A952AD5AB54A952AD5AA54A956AD5AB54A952AD5AB56A952A54AB56AD5AB54A952A54AB56AD5AB54A952A54A952AD5AB56AD5AB56A952A54A952A54A952AD5AB56AD5AB56AD5AB56A952A54A952A54A952A54A952A54";

cyclonev_ram_block ram_block1a128(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a128_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a128.clk0_core_clock_enable = "ena0";
defparam ram_block1a128.clk0_input_clock_enable = "ena0";
defparam ram_block1a128.clk0_output_clock_enable = "ena0";
defparam ram_block1a128.data_interleave_offset_in_bits = 1;
defparam ram_block1a128.data_interleave_width_in_bits = 1;
defparam ram_block1a128.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a128.init_file_layout = "port_a";
defparam ram_block1a128.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a128.operation_mode = "rom";
defparam ram_block1a128.port_a_address_clear = "none";
defparam ram_block1a128.port_a_address_width = 13;
defparam ram_block1a128.port_a_data_out_clear = "none";
defparam ram_block1a128.port_a_data_out_clock = "clock0";
defparam ram_block1a128.port_a_data_width = 1;
defparam ram_block1a128.port_a_first_address = 40960;
defparam ram_block1a128.port_a_first_bit_number = 8;
defparam ram_block1a128.port_a_last_address = 49151;
defparam ram_block1a128.port_a_logical_ram_depth = 65536;
defparam ram_block1a128.port_a_logical_ram_width = 24;
defparam ram_block1a128.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a128.ram_block_type = "auto";
defparam ram_block1a128.mem_init3 = "000000000000000000007FFFFFFFE0000007FFFFC00003FFFE0001FFFC000FFF8003FFC007FF001FF801FF801FF007FC03FE01FE01FE03FC07F00FE03F01FC0FE07F03F03F03F03F07E07C0F81F07E0F83E07C1F0F83E0F87C1E0F07C3C1E0F0F8787C3C3C3E1E1E1E1E3C3C3C387870F1E1C3C78F0E1C3871E3C70E1C78E3C71E38E1C71C38E38E38E38E38E38E38E31C71C638E71C638C738E718E718E718C739CE318C6318C6318C6339CE6319CE63398CE63399CC663399CCC66333998CCC666733319999CCCCCCC66666666666666666666666664CCCCCC9999933326664CCD99B33666CC99B3264CD9B366CD9B366C99326C99364D9B26C9B26D9364DB";
defparam ram_block1a128.mem_init2 = "26D936C936C936C936D924DB6C9249B6DB6492492492492492492492DB6DB4924B6DA492DB492DA496D25B496D25A4B696D2D25A5B4B4B4B496969694B4B4B4A5A5AD2D694B4A52D694A5AD6B4A5294A5294A56B5A94A56B5295A95AD4AD4AD4A95A952B56A54A952A54A956AD52AD5AA552AD52A954AA552AB552AB552AA554AAB554AAA5552AAB5552AAAD5556AAAAD55556AAAAA95555555AAAAAAAAAAB555555555555555555555555555556AAAAAAAAAAD5555554AAAAAB55555AAAAB5555AAAA5554AAAD556AAB554AA9556AAD54AAD54AAD56AB55AAD56A956A956A956AD52A54A952A54A952B56A56AD4AD4AD4AD4AD6A56B5295AD4A5295AD6B5AD6";
defparam ram_block1a128.mem_init1 = "B5AD294A52D6B4A5AD296B4B5A5AD2D296969694B4B4B4B6969696D2D2DA5B4B696D2DA4B692DA4B6925B492DB4925B6D2496DB6D24924925B6DB6DB6DB6D924924936DB6C924DB6C926DB24DB649B649B24D926C9364D926C9B26C9B364D9326C99366CD93264C993264CD9B3266CC99B33664CCD99B3326664CCCD9999B33333266666666666666666666666666666733333319999CCCCE6663331998CCE6633198CC6633198CE63399CC63398CE7318CE7318C6339CE739CE739C6318C739C631CE31CE31CE31C639C738E31C738E39C71C718E38E38E38E38E38E38E1C71C70E38F1C70E3871E3871E3870E3C78F1E3C78F0E1C3C7870F1E1E1C3C3C7878";
defparam ram_block1a128.mem_init0 = "7878787878787C3C3C1E1E0F0F87C3C1E0F07C3E0F07C3E0F83E0F83E0F83E0FC1F07E0FC1F83F03E07E07E07E07E07E07F03F81FC07E03F80FE03FC07F00FF01FE01FE00FF007F803FE007FC00FFC00FFC007FF001FFE001FFE000FFFC000FFFE0003FFFE00007FFFF000003FFFFFC0000001FFFFFFFFF00000000000000001FFFFFFFFFFFFFFF00000000000000001FFFFFFFFF80000007FFFFFC00000FFFFF00003FFFE0001FFFC000FFFC001FFF000FFF001FFE007FF003FF003FF007FE00FF803FC01FE01FF00FE01FE03FC07F80FE03F80FE03F01FC0FE07E03F03F03F03F03F03E07E07C0F81F03E0FC1F07E0F83E0F83E0F83E0F07C1F0F83C1E0F87";

cyclonev_ram_block ram_block1a152(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a152_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a152.clk0_core_clock_enable = "ena0";
defparam ram_block1a152.clk0_input_clock_enable = "ena0";
defparam ram_block1a152.clk0_output_clock_enable = "ena0";
defparam ram_block1a152.data_interleave_offset_in_bits = 1;
defparam ram_block1a152.data_interleave_width_in_bits = 1;
defparam ram_block1a152.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a152.init_file_layout = "port_a";
defparam ram_block1a152.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a152.operation_mode = "rom";
defparam ram_block1a152.port_a_address_clear = "none";
defparam ram_block1a152.port_a_address_width = 13;
defparam ram_block1a152.port_a_data_out_clear = "none";
defparam ram_block1a152.port_a_data_out_clock = "clock0";
defparam ram_block1a152.port_a_data_width = 1;
defparam ram_block1a152.port_a_first_address = 49152;
defparam ram_block1a152.port_a_first_bit_number = 8;
defparam ram_block1a152.port_a_last_address = 57343;
defparam ram_block1a152.port_a_logical_ram_depth = 65536;
defparam ram_block1a152.port_a_logical_ram_width = 24;
defparam ram_block1a152.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a152.ram_block_type = "auto";
defparam ram_block1a152.mem_init3 = "C3E0F0783E1F07C1E0F83E0F83E0F83E0FC1F07E0F81F03E07C0FC0F81F81F81F81F81F80FC0FE07F01F80FE03F80FE03FC07F80FF00FE01FF00FF007F803FE00FFC01FF801FF801FFC00FFF001FFE001FFF0007FFE0007FFF0000FFFF80001FFFFE000007FFFFFC0000003FFFFFFFFF00000000000000001FFFFFFFFFFFFFFF00000000000000001FFFFFFFFF00000007FFFFF800001FFFFC0000FFFF8000FFFE0007FFE000FFF000FFF001FFC007FE007FE007FC00FF803FC01FE00FF00FF01FE01FC07F80FE03F80FC07F03F81FC0FC0FC0FC0FC0FC0F81F83F07E0FC1F07E0F83E0F83E0F83E0F87C1E0F87C1E0F0787C3E1E0F0F078787C3C3C3C3C3C3C";
defparam ram_block1a152.mem_init2 = "3C3C787870F0F1E1C3C7870E1E3C78F1E3C78E1C38F1C38F1C38E1C71E38E1C71C70E38E38E38E38E38E38E31C71C738E39C718E39C738C718E718E718E718C739C6318C739CE739CE7398C6319CE6319CE63398C673398CE633198CC6633198CCE663331998CCCE666733331999999CCCCCCCCCCCCCCCCCCCCCCCCCCCCCC999999B333366664CCC999B336664CD99B3266CC99B3664C993264C99366CD9326C99364D9B26C9B26C9364D926C93649B24DB24DB649B6C926DB64926DB6D924924936DB6DB6DB6DB492492496DB6D2496DB4925B6925B492DA4B692DA4B696D2DA5B4B69696D2D2D2DA5A5A5A52D2D2D29696B4B5A5AD296B4A5AD694A5296B5A";
defparam ram_block1a152.mem_init1 = "D6B5AD6B5294A56B5295AD4AD6A56A56A56A56AD4AD5A952A54A952A54A956AD52AD52AD52AD56AB55AAD56AA556AA556AAD552AA555AAAD556AAA5554AAAB5555AAAAB55555AAAAAA55555556AAAAAAAAAAD55555555555555555555555555555AAAAAAAAAAB55555552AAAAAD55556AAAAD5556AAA9555AAA9554AAA555AAA554AA955AA955AA954AA552A956A954AB56A956AD52A54A952A54AD5A952B52A56A56A56B52B5295AD4A52B5AD4A5294A5294A5AD6B4A52D694A5A52D696B4B4A5A5A5A52D2D2D25A5A5A5B4B49696D2DA4B496D25B496D24B6925B6924B6DA4925B6DB6924924924924924924924DB6DB24926DB64936D926D926D926D936C9";
defparam ram_block1a152.mem_init0 = "B64D936C9B26C9B364D9326C99326CD9B366CD9B3664C99B3266CCD99B336664CCC9999333326666664CCCCCCCCCCCCCCCCCCCCCCCCC666666733331999CCCC666333998CC6673398CC673398CE63398CE7318CE7398C6318C6318C6318E739C631CE31CE31CE39C638C71CE38C71C718E38E38E38E38E38E38E3871C70E38F1C78E3C70E1C78F1C3870E1E3C7870F1E1C3C38787878F0F0F0F0F878787C3C3E1E0F0787C1E0F07C3E0F83E1F07C0F83E0FC1F03E07C0FC1F81F81F81F81FC0FE07F01F80FE01FC07F80FF00FF00FF807FC01FF003FF003FF001FFC007FF8003FFE0007FFF0000FFFF800007FFFFC000000FFFFFFFFC00000000000000000000";

cyclonev_ram_block ram_block1a176(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a176_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a176.clk0_core_clock_enable = "ena0";
defparam ram_block1a176.clk0_input_clock_enable = "ena0";
defparam ram_block1a176.clk0_output_clock_enable = "ena0";
defparam ram_block1a176.data_interleave_offset_in_bits = 1;
defparam ram_block1a176.data_interleave_width_in_bits = 1;
defparam ram_block1a176.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a176.init_file_layout = "port_a";
defparam ram_block1a176.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a176.operation_mode = "rom";
defparam ram_block1a176.port_a_address_clear = "none";
defparam ram_block1a176.port_a_address_width = 13;
defparam ram_block1a176.port_a_data_out_clear = "none";
defparam ram_block1a176.port_a_data_out_clock = "clock0";
defparam ram_block1a176.port_a_data_width = 1;
defparam ram_block1a176.port_a_first_address = 57344;
defparam ram_block1a176.port_a_first_bit_number = 8;
defparam ram_block1a176.port_a_last_address = 65535;
defparam ram_block1a176.port_a_logical_ram_depth = 65536;
defparam ram_block1a176.port_a_logical_ram_width = 24;
defparam ram_block1a176.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a176.ram_block_type = "auto";
defparam ram_block1a176.mem_init3 = "54A952A54A952A54A952A54A952AD5AB56AD5AB56AD5AB56A952A54A952A54A952AD5AB56AD5AB56A952A54A952A55AB56AD5AA54A952A55AB56AD5AA54A952AD5AB56A952A55AB56AD52A54AB56A952A55AB56A952AD5AB54A956AD52A55AB54A956AD52AD5AA54AB56A956AD52AD5AA55AA54AB54A956A956A956AD52AD52AD52AD52AD52AD52AD52AD52AD52AD52AD56A956A954AB54AB55AA552AD52A956AB54AA55AAD52A954AB55AAD56A954AA552A954AA552A954AA552A954AA556AB55AA954AA556AB552A955AA954AAD54AAD54AAD54AAD54AAD54AAD55AA955AAB552AA556AAD55AAB556AAD55AAB556AAD552AA555AAB554AAB556AA9554AAB55";
defparam ram_block1a176.mem_init2 = "4AAB555AAAD552AA9554AAA5556AAB5552AA9555AAA95552AAB5556AAAD555AAAB5554AAA95554AAAB5555AAAAD5556AAAA55556AAAAD5555AAAAB55554AAAAA555556AAAAA555554AAAAAB555555AAAAAAB5555554AAAAAAAD55555552AAAAAAAAD555555555AAAAAAAAAAAB555555555555552AAAAAAAAAAAAAAAAAAAAAAD555555555555555555555555555555555555552AAAAAAAAAAAAAAAAAAAAA955555555555556AAAAAAAAAA9555555554AAAAAAAAD5555554AAAAAA9555555AAAAAA555554AAAAAD55556AAAA955552AAAB55552AAA95554AAAB5554AAA95552AAA5556AAA5556AAA5552AA9556AAB554AAB554AAB556AA9552AA554AA955AAB552";
defparam ram_block1a176.mem_init1 = "AB552AB552AB552A955AAD56AB552A956AB55AAD52A956AB54AB54AB54AB54AB54AB56A952AD5AA54AB56AD5AB56AD5AB56AD5AB56A54A95AB52A56AD4AD5A95A952B52B52B52B52B52B52B5A95A94AD4A56A52B5A94AD6B5295AD6B5294A56B5AD6B5AD6B5AD6B5AD6B5AD6B4A5296B5AD294B5AD296B4A52D694B4A5AD29694B4A5A52D2D69696B4B4B4A5A5A5A5A5A5A5A5A5A5A5A5A5A4B4B4B6969692D2DA5A4B49692D25A4B696D25A4B692DA4B692DA4B6D25B692DB492DA496DB492DB6924B6DA4925B6DB492496DB6DB6D24924924924924924924924924924DB6DB6D924924DB6D9249B6D9249B6C926DB249B649B6C936C936C93649B64DB26D93";
defparam ram_block1a176.mem_init0 = "649B26C9364D9364D9364D9364D9326C9B364D9B264D9B264C9B366CD9B366CD9B3664C99B3664CD9B32664CD99332664CC9993336664CCD999B33326666CCCCC999999B3333333366666666666666666666666666666666333333333999998CCCCC666673331999CCCE667333998CCE6633198CCE673398CC663398CC67319CC67319CE6339CC6339CC6319CE7398C6318C6318C6318E739CE318C739C639CE31CE31CE31CE39C638C718E39C718E39C71CE38E39C71C71C71CE38E38E38E1C71C71C71E38E3871C70E38F1C78E1C70E3C70E3C78E1C3870E1C3870E1C3C78F0E1E3C387870F0E1E1E1E3C3C3C3C3C3C3C3C3C1E1E1E0F0F0787C3C1E0F0F87";

cyclonev_ram_block ram_block1a56(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a56_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a56.clk0_core_clock_enable = "ena0";
defparam ram_block1a56.clk0_input_clock_enable = "ena0";
defparam ram_block1a56.clk0_output_clock_enable = "ena0";
defparam ram_block1a56.data_interleave_offset_in_bits = 1;
defparam ram_block1a56.data_interleave_width_in_bits = 1;
defparam ram_block1a56.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a56.init_file_layout = "port_a";
defparam ram_block1a56.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a56.operation_mode = "rom";
defparam ram_block1a56.port_a_address_clear = "none";
defparam ram_block1a56.port_a_address_width = 13;
defparam ram_block1a56.port_a_data_out_clear = "none";
defparam ram_block1a56.port_a_data_out_clock = "clock0";
defparam ram_block1a56.port_a_data_width = 1;
defparam ram_block1a56.port_a_first_address = 16384;
defparam ram_block1a56.port_a_first_bit_number = 8;
defparam ram_block1a56.port_a_last_address = 24575;
defparam ram_block1a56.port_a_logical_ram_depth = 65536;
defparam ram_block1a56.port_a_logical_ram_width = 24;
defparam ram_block1a56.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a56.ram_block_type = "auto";
defparam ram_block1a56.mem_init3 = "3C1F0F87C1E0F83C1F07C1F07C1F07C1F03E0F81F07E0FC1F83F03E07E07E07E07E07E07F03F01F80FE07F01FC07F01FC03F807F00FF01FE00FF00FF807FC01FF007FE007FE007FE003FF000FFE001FFE000FFF8001FFF8000FFFF00007FFFE00001FFFFF8000007FFFFFFC000000000FFFFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFFFE000000000FFFFFFF8000007FFFFE00003FFFF00007FFF0001FFF8001FFF000FFF000FFE003FF801FF801FF803FF007FC03FE01FF00FF00FE01FE03F807F01FC07F03F80FC07E03F03F03F03F03F03F07E07C0F81F03E0F81F07C1F07C1F07C1F0783E1F0783E1F0F8783C1E1F0F0F878783C3C3C3C3C3C3";
defparam ram_block1a56.mem_init2 = "C3C38787870F0E1E3C3878F1E1C3870E1C3871E3C70E3C70E3C71E38E1C71E38E38F1C71C71C71C71C71C71CE38E38C71C638E71C638C738E718E718E718E738C639CE738C6318C6318C6739CE6319CE6319CC63398CC67319CCE673399CCE6733199CCCE66733319998CCCCE6666673333333333333333333333333333336666664CCCC9999B3336664CCD99B32664CD9933664C99B366CD9B366C99326CD9366C9B264D9364D936C9B26D936C9B64DB24DB249B64936D9249B6D924936DB6DB6C92492492492496DB6DB692492DB6924B6DA496DA4B6D25B496D25B49692DA5A4B49696D2D2D2D25A5A5A5A52D2D2D69694B4A5A52D694B5A5296B5AD694A5";
defparam ram_block1a56.mem_init1 = "294A5294AD6B5A94AD6A52B5295A95A95A95A952B52A56AD5AB56AD5AB56A952AD52AD52AD52A954AA552A955AA955AA9552AAD55AAA5552AA9555AAAB5554AAAA55554AAAAA555555AAAAAAA955555555552AAAAAAAAAAAAAAAAAAAAAAAAAAAAA55555555554AAAAAAAD555552AAAA955552AAA95556AAA5556AAA555AAA555AAB556AA556AA556AB55AAD56A956AB54A956A952AD5AB56AD5AB52A56AD4AD5A95A95A94AD4AD6A52B5AD4A52B5AD6B5AD6B5A5294B5AD296B5A5AD29694B4B5A5A5A5AD2D2D2D25A5A5A4B4B69692D25B4B692DA4B692DB496DA496DB4925B6DA4924B6DB6DB6DB6DB6DB6DB6DB24924DB6D9249B6C926D926D926D926C936";
defparam ram_block1a56.mem_init0 = "49B26C9364D9364C9B26CD9366C993264C993264C99B3664CD99332664CC999B3336666CCCCD999999B33333333333333333333333339999998CCCCE6663333999CCC66733998CC673399CC67319CC67318CE7318C6739CE739CE739CE718C639CE31CE31CE31CE39C738E31C738E38E71C71C71C71C71C71C71C78E38F1C70E3871C38F1E3870E3C78F1E1C3878F1E1E3C3C78787870F0F0F0F07878787C3C1E1F0F8783E1F0F83C1F07C1E0F83F07C1F03E0FC1F83F07E07E07E07E07E03F01F80FE07F01FE03F807F00FF00FF007F803FE00FFC00FFC00FFE003FF8007FFC001FFF8000FFFF00007FFFF800003FFFFFF000000003FFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a80(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a80_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a80.clk0_core_clock_enable = "ena0";
defparam ram_block1a80.clk0_input_clock_enable = "ena0";
defparam ram_block1a80.clk0_output_clock_enable = "ena0";
defparam ram_block1a80.data_interleave_offset_in_bits = 1;
defparam ram_block1a80.data_interleave_width_in_bits = 1;
defparam ram_block1a80.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a80.init_file_layout = "port_a";
defparam ram_block1a80.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a80.operation_mode = "rom";
defparam ram_block1a80.port_a_address_clear = "none";
defparam ram_block1a80.port_a_address_width = 13;
defparam ram_block1a80.port_a_data_out_clear = "none";
defparam ram_block1a80.port_a_data_out_clock = "clock0";
defparam ram_block1a80.port_a_data_width = 1;
defparam ram_block1a80.port_a_first_address = 24576;
defparam ram_block1a80.port_a_first_bit_number = 8;
defparam ram_block1a80.port_a_last_address = 32767;
defparam ram_block1a80.port_a_logical_ram_depth = 65536;
defparam ram_block1a80.port_a_logical_ram_width = 24;
defparam ram_block1a80.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a80.ram_block_type = "auto";
defparam ram_block1a80.mem_init3 = "AB56AD5AB56AD5AB56AD5AB56AD52A54A952A54A952A54A956AD5AB56AD5AB56AD52A54A952A54A956AD5AB56AD5AA54A952A54AB56AD5AB54A952A55AB56AD52A54A956AD5AA54A952AD5AB54A952AD5AA54A956AD52A54AB56A952AD5AA54AB56A952AD5AA55AB54A956A952AD52A55AA54AB54AB56A956A956AD52AD52AD52AD52AD52AD52AD52AD52AD52AD52AD52A956A956AB54AB54AA55AA552AD56A954AB55AA552AD56AB54AA552A956AB55AAD56AB55AAD56AB55AAD56AB55AA954AA556AB55AA954AAD56AA556AB552AB552AB552AB552AB552AB552AB556AA554AAD55AA9552AA554AA9552AA554AA9552AAD55AAB554AAB554AA9556AA9554AA";
defparam ram_block1a80.mem_init2 = "B554AAA555AAAD556AAB555AAA9554AAAD556AAA5556AAAD554AAA95552AAA5554AAAB5556AAAB5554AAAA55552AAA95555AAAA95555AAAAA55554AAAAB55555AAAAAD55555AAAAAB555554AAAAAA5555554AAAAAAB55555552AAAAAAAD555555552AAAAAAAAA555555555554AAAAAAAAAAAAAAD5555555555555555555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAD5555555555555555555556AAAAAAAAAAAAA955555555556AAAAAAAAB555555552AAAAAAB5555556AAAAAA555555AAAAAB555552AAAA955556AAAAD5554AAAAD5556AAAB5554AAAB5556AAAD555AAA9555AAA9555AAAD556AAB554AAB554AAB554AA9556AAD55AAB556AA554AAD";
defparam ram_block1a80.mem_init1 = "54AAD54AAD54AAD56AA552A954AAD56A954AA552AD56A954AB54AB54AB54AB54AB54A956AD52A55AB54A952A54A952A54A952A54A95AB56A54AD5A952B52A56A54AD4AD4AD4AD4AD4AD4AD4A56A56B52B5A95AD4A56B5294AD6A5294AD6B5A94A5294A5295AD694A5294A5294B5AD694A52D6B4A52D694B5AD296B4B5A52D696B4B5A5AD2D2969694B4B4B5A5A5A5A5A5A5A5A5A5A5A5A5A5B4B4B4B69696D2D25A5B4B696D2DA5B49692DA5B496D25B496D25B492DA496D24B6925B6924B6D2496DB4925B6DA4924B6DB692492496DB6DB6DB6DB6DB6DB6DB6DB6DB6DB64924926DB6DB24926DB64926DB64936D924DB649B64936C936C936C9B649B24D926C";
defparam ram_block1a80.mem_init0 = "9B64D936C9B26C9B26C9B26C9B26CD9364C9B264D9B264D9B364C993264C993264C99B3664C99B3264CD99B3266CCD99B33666CCC999B3326664CCCD9999333336666664CCCCCCCD99999999999999999999999999999999CCCCCCCCC6666663333399998CCCE6663331998CCC66733199CCE6733198CC673399CC673398CE63398CE6319CC6339CC6339CE6318C6739CE739CE739CE718C631CE738C639C631CE31CE31CE31C639C738E71C638C71C638E31C71C638E38E38E71C71C71C71C38E38E38E1C71C78E38F1C70E3871E38F1C38F1C3871E3C78F1E3C78F1E3C3870F1E1C3C7878F0F1E1E1E1C3C3C3C3C3C3C3C3C3E1E1E1F0F0F8783C3E1E0F078";

cyclonev_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "rom";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "clock0";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 8191;
defparam ram_block1a8.port_a_logical_ram_depth = 65536;
defparam ram_block1a8.port_a_logical_ram_width = 24;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init3 = "3C1E0F0F8783C3E1E1F0F0F0F8787878787878787870F0F0F1E1E3C3C7870F1E1C3878F1E3C78F1E3C78F1C3871E3871E38F1C38E1C71E38E3C71C70E38E38E3871C71C71C71CE38E38E38C71C718E38C71C638C71CE39C738C718E718E718E718C738C639CE718C631CE739CE739CE739CC6318CE7398C67398C67318CE63398CE63399CC673399CC6633199CCE6733199CCC6663331998CCCE6663333399998CCCCCC66666666733333333333333333333333333333333666666664CCCCCD99999333366664CCC999B332666CCD99B33666CC99B33664C99B3264CD9B3264C993264C993264D9B364C9B364C9B264D9366C9B26C9B26C9B26C9B26D9364DB2";
defparam ram_block1a8.mem_init2 = "6C93649B24DB26D926D926D924DB24DB64936D924DB6C924DB6C9249B6DB6C924924DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6D2492492DB6DA4924B6DB4925B6D2496DA492DB492DA496D24B6925B496D25B496D25B4B692D25B4B696D2DA5B4B49696D2D2DA5A5A5B4B4B4B4B4B4B4B4B4B4B4B4B4B5A5A5A52D2D29696B4B5A5AD2D694B5A5AD296B5A52D694A5AD694A52D6B5A5294A5294A52D6B5294A5294A52B5AD6A5294AD6A5295AD4A56B52B5A95AD4AD4A56A56A56A56A56A56A56A54AD4A95A952B56A54AD5AB52A54A952A54A952A54A952A55AB54A956AD52A55AA55AA55AA55AA55AA552AD56A954AA552AD56AA552A954AAD56AA556AA556AA55";
defparam ram_block1a8.mem_init1 = "6AA554AAD55AAB556AAD552AA555AAA555AAA555AAAD556AAB5552AAB5552AAB5556AAAD555AAAA5555AAAAD5556AAAA55556AAAAD55552AAAA955555AAAAAB555554AAAAAAD555555AAAAAAA955555555AAAAAAAAAD55555555552AAAAAAAAAAAAAD5555555555555555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAB55555555555555555555556AAAAAAAAAAAAAA555555555554AAAAAAAAA9555555556AAAAAAA95555555AAAAAAA5555554AAAAAA555555AAAAAB555556AAAAB55555AAAAA55554AAAAB55552AAAB55552AAA95554AAAA5555AAAAD555AAAA5554AAA95552AAA5556AAAD554AAAD556AAA5552AAB555AAAD556AAB554AAA555A";
defparam ram_block1a8.mem_init0 = "AA5552AAD552AA555AAA555AAB556AA9552AA554AA9552AA554AA9552AB556AA554AAD55AA955AA955AA955AA955AA955AA955AAD54AAD56AA552AB55AAD54AA552AB55AAD56AB55AAD56AB55AAD56AB55AAD52A954AA55AAD56A954AB55AA552AD56A954AB54AA55AA55AAD52AD52A956A956A956A956A956A956A956A956A956A956A956AD52AD52AD5AA55AA54AB54A956A952AD52A55AB54AB56A952AD5AA54AB56A952AD5AA54A956AD52A54AB56A952A55AB56A952A54AB56AD52A54A956AD5AB54A952A55AB56AD5AA54A952A54AB56AD5AB56AD52A54A952A54A956AD5AB56AD5AB56AD52A54A952A54A952A54A956AD5AB56AD5AB56AD5AB56AD5AA";

cyclonev_ram_block ram_block1a32(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a32_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a32.clk0_core_clock_enable = "ena0";
defparam ram_block1a32.clk0_input_clock_enable = "ena0";
defparam ram_block1a32.clk0_output_clock_enable = "ena0";
defparam ram_block1a32.data_interleave_offset_in_bits = 1;
defparam ram_block1a32.data_interleave_width_in_bits = 1;
defparam ram_block1a32.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a32.init_file_layout = "port_a";
defparam ram_block1a32.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a32.operation_mode = "rom";
defparam ram_block1a32.port_a_address_clear = "none";
defparam ram_block1a32.port_a_address_width = 13;
defparam ram_block1a32.port_a_data_out_clear = "none";
defparam ram_block1a32.port_a_data_out_clock = "clock0";
defparam ram_block1a32.port_a_data_width = 1;
defparam ram_block1a32.port_a_first_address = 8192;
defparam ram_block1a32.port_a_first_bit_number = 8;
defparam ram_block1a32.port_a_last_address = 16383;
defparam ram_block1a32.port_a_logical_ram_depth = 65536;
defparam ram_block1a32.port_a_logical_ram_width = 24;
defparam ram_block1a32.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.ram_block_type = "auto";
defparam ram_block1a32.mem_init3 = "FFFFFFFFFFFFFFFFFFFF800000001FFFFFF800003FFFFC0001FFFE0003FFF0007FFC003FF800FFE007FE007FE00FF803FC01FE01FE01FC03F80FF01FC0FE03F01F80FC0FC0FC0FC0FC1F83F07E0F81F07C1F83E0F07C1F0783E1F0F83C3E1F0F0787C3C3C3C1E1E1E1E1C3C3C3C7878F0F1E3C3870F1E3C78E1C38F1E3871C38E1C71E38E3C71C71C71C71C71C71C71CE38E39C718E39C738E718E718E718E738C631CE739CE739CE739CC6319CE6319CC67319CC673399CC6633399CCC6673339998CCCE666633333339999999999999999999999999B33333366666CCCD999B332664CC99933664CD9B3264C993264C99326CD9366C9B264D9364D926C9B24";
defparam ram_block1a32.mem_init2 = "D926C936C936C936C926DB24936DB649249B6DB6DB6DB6DB6DB6DB6DA4924B6DB4925B6D24B6D25B692DA4B692DA5B49692D2DA5A4B4B4B496969696B4B4B4B5A5A52D296B4B5AD296B5A5294B5AD6B5AD6B5A94A56B5A94AD6A56A52B52B52B56A56AD4A95AB56AD5AB56A952AD52A55AAD52AD56AB55AAD54AAD54AAD55AAB554AAB554AAAD554AAAD5552AAA955552AAAA9555556AAAAAAA55555555554AAAAAAAAAAAAAAAAAAAAAAAAAAAAA955555555552AAAAAAB555554AAAAA55554AAAA5555AAAB5552AA9554AAB556AA9552AB552AB552A954AA552A956A956A956A952AD5AB56AD5AB56AD4A95A952B52B52B52B5295A94AD6A52B5AD6A5294A529";
defparam ram_block1a32.mem_init1 = "4A52D6B5AD294B5A52D694B4A5A52D2D6969694B4B4B4B496969696D2D25A4B4B692D25B496D25B496DA4B6D24B6DA492DB692492DB6DB6D24924924924926DB6DB6D924936DB24936D924DB249B649B64DB26D936C9B26D9364D9364C9B26CD9366C99326CD9B366CD9B3264CD9933664CC99B336664CCD999B333266664CCCCCD999999999999999999999999999999CCCCCCE666633331999CCCE66733199CCE673399CCE67319CC663398C67318CE7318CE739CC6318C6318C639CE738C639CE31CE31CE31CE39C638C71CE38C71C638E38E71C71C71C71C71C71C71E38E38F1C70E38F1C78E1C78E1C78F1C3870E1C3870F1E3C3878F0E1E1C3C3C38787";
defparam ram_block1a32.mem_init0 = "87878787878783C3C3E1E1F0F0783C3E1F0F83C1F0F83C1F07C1F07C1F07C1F03E0F81F03E07C0FC1F81F81F81F81F81F80FC07E03F81FC07F01FC03F80FF00FE01FE01FF00FF807FC01FF803FF003FF003FF800FFE001FFE001FFF0003FFF0001FFFC0001FFFF80000FFFFFC000003FFFFFFE000000000FFFFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFFFE0000000007FFFFFFC000003FFFFF00000FFFFC0001FFFE0003FFF0003FFE000FFF000FFE001FF800FFC00FFC00FFC01FF007FC03FE01FE00FF01FE01FC03F807F01FC07F01FC0FE03F01F81FC0FC0FC0FC0FC0FC0F81F83F07E0FC1F03E0F81F07C1F07C1F07C1F0783E0F07C3E1F078";

cyclonev_ram_block ram_block1a105(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a105_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a105.clk0_core_clock_enable = "ena0";
defparam ram_block1a105.clk0_input_clock_enable = "ena0";
defparam ram_block1a105.clk0_output_clock_enable = "ena0";
defparam ram_block1a105.data_interleave_offset_in_bits = 1;
defparam ram_block1a105.data_interleave_width_in_bits = 1;
defparam ram_block1a105.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a105.init_file_layout = "port_a";
defparam ram_block1a105.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a105.operation_mode = "rom";
defparam ram_block1a105.port_a_address_clear = "none";
defparam ram_block1a105.port_a_address_width = 13;
defparam ram_block1a105.port_a_data_out_clear = "none";
defparam ram_block1a105.port_a_data_out_clock = "clock0";
defparam ram_block1a105.port_a_data_width = 1;
defparam ram_block1a105.port_a_first_address = 32768;
defparam ram_block1a105.port_a_first_bit_number = 9;
defparam ram_block1a105.port_a_last_address = 40959;
defparam ram_block1a105.port_a_logical_ram_depth = 65536;
defparam ram_block1a105.port_a_logical_ram_width = 24;
defparam ram_block1a105.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a105.ram_block_type = "auto";
defparam ram_block1a105.mem_init3 = "954AB55AAD56A954AB55AA55AAD52AD52AD52AD52AD5AA55AB54A956AD52A54AB56AD5AB56AD5AB56AD5AB56AD4A952B56A54A95AB52B56A56AD4AD5A95A95A95AB52B52B52B5A95A95A95AD4AD4A56A52B5A95AD4A56B5295AD4A52B5AD4A52B5AD6A5294A52B5AD6B5AD6B5AD6B5AD6B5AD6B5A5294A52D6B5AD294A5AD694A5AD694B5AD296B4A52D694B4A5AD296B4B5A52D29694B4A5A5AD2D69696B4B4B5A5A5AD2D2D2D2D696969696969696969696969696969692D2D2D2D25A5A5B4B4B49696D2D2DA5A4B49696D2DA5B4B696D2DA5B49692D25B49692DA4B696D25B496D25B496D24B692DA496D25B692DB492DA496DA496DA496DA496DB492DB69";
defparam ram_block1a105.mem_init2 = "25B6D2496DB6924B6DB4924B6DB692492DB6DB4924925B6DB6DA4924924925B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB64924924926DB6DB6C924924DB6DB64924DB6DB24926DB6C924DB6C924DB6C926DB64936D924DB64936D924DB249B64936C936D926D926D926D926D926D926D936C936C9B649B24D926C93649B24D936C9B64D936C9B24D9364DB26C9B26C9364D9364D9364D9364D9364D9366C9B26C9B264D9364C9B26CD9366C9B364D9B26CD9326CD9326CD9326CD9B264D9B364C99326CD9B366C993264C993264C993264C993366CD9B3264C993366CC993366CC993366CC99B3264CD9933664CD9933664CD99B3266CCD9933266CC";
defparam ram_block1a105.mem_init1 = "D99332664CC999332664CC999333666CCC9993336664CCD9993336666CCC999933326664CCC9999333366664CCCD99993333266664CCCC99999B33333666666CCCCCD999999B33333366666664CCCCCCCC999999999B3333333333666666666666664CCCCCCCCCCCCCCCCCCCCCD999999999999999999999999999999999999998CCCCCCCCCCCCCCCCCCCCCCE666666666666663333333333339999999998CCCCCCCCE6666666733333339999999CCCCCCC666666333333999998CCCCCE666673333399999CCCCC66667333319998CCCCE666733339999CCCC666633339999CCCC66673331999CCCE6663333999CCCE6663331998CCC6663331998CCC6663339";
defparam ram_block1a105.mem_init0 = "99CCC666333199CCC666333998CCE66733199CCC66733199CCC66733198CCE6633399CCC66733998CC66733998CC66733998CC6633399CCE6633198CC6633399CCE673399CCE673399CCE673399CCE673399CCE673399CC6633198CC673399CCE633198CE673399CC663399CCE633198CE673198CE673198CE673198CE673198CE673198CE63319CCE63399CC673398CC673198CE63319CC673398CE67319CC663398CE67319CC663398CE63319CC67319CCE63398CE67319CC67319CCE63398CE63398CC67319CC67319CC673398CE63398CE63398CE63319CC67319CC67319CC67319CC67319CCE63398CE63398CE63398CE63398CE63398CE63398CE63398";

cyclonev_ram_block ram_block1a129(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a129_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a129.clk0_core_clock_enable = "ena0";
defparam ram_block1a129.clk0_input_clock_enable = "ena0";
defparam ram_block1a129.clk0_output_clock_enable = "ena0";
defparam ram_block1a129.data_interleave_offset_in_bits = 1;
defparam ram_block1a129.data_interleave_width_in_bits = 1;
defparam ram_block1a129.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a129.init_file_layout = "port_a";
defparam ram_block1a129.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a129.operation_mode = "rom";
defparam ram_block1a129.port_a_address_clear = "none";
defparam ram_block1a129.port_a_address_width = 13;
defparam ram_block1a129.port_a_data_out_clear = "none";
defparam ram_block1a129.port_a_data_out_clock = "clock0";
defparam ram_block1a129.port_a_data_width = 1;
defparam ram_block1a129.port_a_first_address = 40960;
defparam ram_block1a129.port_a_first_bit_number = 9;
defparam ram_block1a129.port_a_last_address = 49151;
defparam ram_block1a129.port_a_logical_ram_depth = 65536;
defparam ram_block1a129.port_a_logical_ram_width = 24;
defparam ram_block1a129.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a129.ram_block_type = "auto";
defparam ram_block1a129.mem_init3 = "00000000000000000000000000001FFFFFFFFFFFC000000001FFFFFFFC0000007FFFFFC00000FFFFF800007FFFF00003FFFE0001FFFE0003FFF0001FFF0003FFE000FFF000FFF000FFE003FF800FFE007FE003FF007FE007FC01FF003FC01FF007F803FC03FE01FE01FE03FC03F807F00FE03FC07F01FC07F01FC0FE03F81FC0FE07E03F03F81F81F81F81F81F81F81F03F03E07E0FC1F83F07E0F81F07E0F83F07C1F07C1F07C1F07C1F07C1E0F83E1F0783E1F0783C1E0F87C3C1E0F0787C3C1E1F0F0F8787C3C3C3C1E1E1E1E1E1E1E1E1E1E1E1E1C3C3C3C787870F0E1E1C3C3878F0E1E3C7870E1C3C78F1E3C78F1E3870E1C78F1C3871E3871E38F1C38";
defparam ram_block1a129.mem_init2 = "E1C70E38F1C70E38F1C71C38E38E3871C71C71C71C71C71C71C71C71C71C738E38E39C71C738E39C71CE38C71CE39C718E31CE39C738C738C718E718C738C739C639CE318C739CE318C639CE739CE739CE739CE7398C6318CE7398C6339CC63398C67318CE63398CE63398CE63319CC663319CCE673399CCE6733198CCE66333998CCC6663331998CCCE666333319999CCCCCE666667333333399999999998CCCCCCCCCCCCCCCCCCCCCCCCCCCCCD9999999999B3333332666666CCCCC9999933336666CCCD999B332666CCD99B332664CD99B32664CD9933664CD9B3264CD9B3264C993264C993264C99326CD9B264D9B264D9B26CD9364C9B26C9B364D9364D";
defparam ram_block1a129.mem_init1 = "93649B26C9B26D93649B26D936C9B649B24DB24D926D926DB24DB249B64936D924DB64926DB64926DB6C9249B6DB6C924924DB6DB6DB6DB6C924924924924B6DB6DB6DB6DA4924925B6DB692492DB6D2496DB4925B6D24B6DA496DA496D24B6925B492DA4B692DA4B692DA4B696D25A4B696D2DA5B4B69692D2DA5A4B4B496969692D2D2D2D2D2D2D2D2D2D2D2D2D2D2D6969694B4B4A5A5AD2D696B4B5A5AD296B4A5AD296B4A5AD694B5AD694A5AD6B5A5294A5296B5AD6B5AD6B5294A5294AD6B5A94A56B5A94AD6B5295A94AD6A56B52B52B5A95A95A95A95A95A95AB52B52A56A54AD5A952B56AD4A952A56AD5AB56AD5AA54A952AD5AB54AB56A952AD5";
defparam ram_block1a129.mem_init0 = "2AD52AD52AD52A956AB54AA55AAD56AB55AAD56AA552A955AA955AA955AA955AAB552AA554AA9556AAD552AAD552AAD552AA9554AAAD556AAA5556AAAD555AAAB5554AAAA55552AAA955552AAAA55555AAAAAD55554AAAAAB555555AAAAAAA55555556AAAAAAAAD5555555556AAAAAAAAAAAAB55555555555555555555555554AAAAAAAAAAAAAAA555555555555555555555555552AAAAAAAAAAAA95555555555AAAAAAAAB55555556AAAAAA9555555AAAAAA555554AAAAA55555AAAAA55554AAAAD5556AAAB5555AAAB5554AAA95552AAB5552AAB555AAA9554AAB555AAA555AAA555AAB554AA9552AA554AA955AAB552AB552AB552AB55AA955AAD56AB552A";

cyclonev_ram_block ram_block1a153(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a153_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a153.clk0_core_clock_enable = "ena0";
defparam ram_block1a153.clk0_input_clock_enable = "ena0";
defparam ram_block1a153.clk0_output_clock_enable = "ena0";
defparam ram_block1a153.data_interleave_offset_in_bits = 1;
defparam ram_block1a153.data_interleave_width_in_bits = 1;
defparam ram_block1a153.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a153.init_file_layout = "port_a";
defparam ram_block1a153.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a153.operation_mode = "rom";
defparam ram_block1a153.port_a_address_clear = "none";
defparam ram_block1a153.port_a_address_width = 13;
defparam ram_block1a153.port_a_data_out_clear = "none";
defparam ram_block1a153.port_a_data_out_clock = "clock0";
defparam ram_block1a153.port_a_data_width = 1;
defparam ram_block1a153.port_a_first_address = 49152;
defparam ram_block1a153.port_a_first_bit_number = 9;
defparam ram_block1a153.port_a_last_address = 57343;
defparam ram_block1a153.port_a_logical_ram_depth = 65536;
defparam ram_block1a153.port_a_logical_ram_width = 24;
defparam ram_block1a153.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a153.ram_block_type = "auto";
defparam ram_block1a153.mem_init3 = "A955AAD56AB552AB55AA955AA955AA955AAB552AA554AA9552AA555AAB554AAB554AAB555AAA5552AAB555AAA9555AAA95552AAA5555AAAB5555AAAAD5556AAAA55554AAAAB55554AAAAA555554AAAAAB5555552AAAAAAD5555555AAAAAAAAB55555555552AAAAAAAAAAAA955555555555555555555555554AAAAAAAAAAAAAAA55555555555555555555555555AAAAAAAAAAAAAD5555555556AAAAAAAAD5555554AAAAAAB555555AAAAAA555556AAAAB55554AAAA955552AAA95554AAAA5555AAAB5556AAAD554AAAD556AAA5552AA9556AA9556AA9556AAD552AA554AA955AAB552AB552AB552AB552A954AAD56AB55AAD56AB54AA55AAD52A956A956A956A9";
defparam ram_block1a153.mem_init2 = "56A952AD5AA55AB56A952A54AB56AD5AB56AD4A952A56AD5A952B56A54AD4A95A95AB52B52B52B52B52B52B5A95A95AD4AD6A52B5295AD6A52B5AD4A52B5AD6A5294A5295AD6B5AD6B5AD294A5294B5AD6B4A52D6B5A52D6B4A5AD296B4A5AD296B4B5A5AD2D696B4B4A5A5A52D2D2D6969696969696969696969696969692D2D2D25A5A4B4B69692D2DA5B4B696D2DA4B496D2DA4B692DA4B692DA4B6925B492DA496D24B6D24B6DA496DB4925B6D2496DB692492DB6DB4924924B6DB6DB6DB6DA4924924924926DB6DB6DB6DB64924926DB6DB24926DB6C924DB6C924DB64936D924DB249B649B6C936C93649B649B24DB26D936C9B24D936C9B26C9B24D93";
defparam ram_block1a153.mem_init1 = "64D9364D9B26C9B264D9366C9B364C9B364C9B366C993264C993264C993264C99B3664C99B3664CD9933664CC99B33664CC999B33666CCC999B3336666CCCD99993333266666CCCCCC9999999B3333333333666666666666666666666666666666333333333339999999CCCCCCE66667333319998CCCE6663331998CCC666333998CCE6633199CCE673399CCE673198CC673198CE63398CE63398CE6319CC63398C67398C6339CE6318C6339CE739CE739CE739CE738C6318E739C6318E738C739C639C631CE31C639C639C738E718E31C738E71C638E71C738E39C71C738E38E39C71C71C71C71C71C71C71C71C71C71C38E38E3871C71E38E1C71E38E1C70E";
defparam ram_block1a153.mem_init0 = "3871E38F1C38F1C3871E3C70E1C38F1E3C78F1E3C7870E1C3C78F0E1E3C387870F0E1E1C3C3C78787870F0F0F0F0F0F0F0F0F0F0F0F07878787C3C3E1E1F0F0787C3C1E0F0787C3E0F0783C1F0F83C1F0F83E0F07C1F07C1F07C1F07C1F07C1F83E0FC1F03E0FC1F83F07E0FC0F81F81F03F03F03F03F03F03F03F81F80FC0FE07F03F80FE07F01FC07F01FC07F80FE01FC03F807F80FF00FF00FF807F803FC01FF007F801FF007FC00FFC01FF800FFC00FFE003FF800FFE001FFE001FFE000FFF8001FFF0001FFF8000FFFF0000FFFF80001FFFFC00003FFFFE000007FFFFFC0000007FFFFFFF0000000007FFFFFFFFFFF00000000000000000000000000000";

cyclonev_ram_block ram_block1a177(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a177_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a177.clk0_core_clock_enable = "ena0";
defparam ram_block1a177.clk0_input_clock_enable = "ena0";
defparam ram_block1a177.clk0_output_clock_enable = "ena0";
defparam ram_block1a177.data_interleave_offset_in_bits = 1;
defparam ram_block1a177.data_interleave_width_in_bits = 1;
defparam ram_block1a177.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a177.init_file_layout = "port_a";
defparam ram_block1a177.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a177.operation_mode = "rom";
defparam ram_block1a177.port_a_address_clear = "none";
defparam ram_block1a177.port_a_address_width = 13;
defparam ram_block1a177.port_a_data_out_clear = "none";
defparam ram_block1a177.port_a_data_out_clock = "clock0";
defparam ram_block1a177.port_a_data_width = 1;
defparam ram_block1a177.port_a_first_address = 57344;
defparam ram_block1a177.port_a_first_bit_number = 9;
defparam ram_block1a177.port_a_last_address = 65535;
defparam ram_block1a177.port_a_logical_ram_depth = 65536;
defparam ram_block1a177.port_a_logical_ram_width = 24;
defparam ram_block1a177.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a177.ram_block_type = "auto";
defparam ram_block1a177.mem_init3 = "3398CE63398CE63398CE63398CE63398CE63398CE63398CE67319CC67319CC67319CC67319CC673198CE63398CE63398CE63399CC67319CC67319CC663398CE63398CE67319CC67319CCE63398CE67319CC673198CE63398CC67319CCE63398CC67319CCE63399CC673198CE63319CC663399CC673398CE673198CE63319CCE63319CCE63319CCE63319CCE63319CCE633198CE673398CC673399CCE633198CE673399CC6633198CC673399CCE673399CCE673399CCE673399CCE673399CCE6733998CC6633198CCE6733998CC6633399CCC6633399CCC6633399CCC66733998CCE6633199CCC66733199CCC66733199CCCE66333998CCC667331998CCC66733";
defparam ram_block1a177.mem_init2 = "3998CCC6663331998CCC6663331998CCCE6673339998CCCE6673331999CCCC666733339998CCCC666733339999CCCCE6666333319999CCCCC666673333399999CCCCCE66666333333999998CCCCCC666666733333339999999CCCCCCCCE666666663333333333999999999998CCCCCCCCCCCCCCE666666666666666666666633333333333333333333333333333333333333366666666666666666666664CCCCCCCCCCCCCD9999999999B333333332666666664CCCCCCD999999B333333666666CCCCCD99999B3333266664CCCC99999333366664CCCD999933326664CCC99993332666CCCD9993336664CCD999332666CCD999332664CC999332664CC999336";
defparam ram_block1a177.mem_init1 = "66CC99933666CC99B33664CD9933664CD9933664C99B3266CD993266CD993266CD993264C99B366CD993264C993264C993264C99326CD9B366C993264D9B364C9B366C99366C99366C99366C9B364D9B26CD9366C9B264D9364C9B26C9B26CD9364D9364D9364D9364D9364D926C9B26C9B64D93649B26D9364DB26D93649B24D926C93649B24DB26D926D936C936C936C936C936C936C936D926D924DB249B64936D924DB64936D924DB6C926DB64926DB64926DB6C9249B6DB64924DB6DB64924926DB6DB6C924924924DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB4924924924B6DB6DB4924925B6DB692492DB6DA4925B6DA492DB6D2496DB49";
defparam ram_block1a177.mem_init0 = "2DB6925B6D24B6D24B6D24B6D24B6925B692DB496D24B692DA496D25B496D25B496D2DA4B692D25B49692D25B4B696D2DA5B4B696D2D25A4B4B69696D2D25A5A5B4B4B49696969692D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D696969696B4B4B5A5A5AD2D2D696B4B4A5A52D29694B5A5AD296B4A5A52D694A5AD296B5A52D6B4A52D6B4A5296B5AD694A5294B5AD6B5AD6B5AD6B5AD6B5AD6B5A94A5294AD6B5A94A56B5A94A56B5295AD4A56B52B5A94AD4A56A56B52B52B52B5A95A95A95AB52B52B52B56A56AD4AD5A95AB52A54AD5A952A56AD5AB56AD5AB56AD5AB56AD5AA54A956AD52A55AB54AB56A956A956A956A956AB54AB55AA552AD56AB55AA552";

cyclonev_ram_block ram_block1a57(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a57_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a57.clk0_core_clock_enable = "ena0";
defparam ram_block1a57.clk0_input_clock_enable = "ena0";
defparam ram_block1a57.clk0_output_clock_enable = "ena0";
defparam ram_block1a57.data_interleave_offset_in_bits = 1;
defparam ram_block1a57.data_interleave_width_in_bits = 1;
defparam ram_block1a57.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a57.init_file_layout = "port_a";
defparam ram_block1a57.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a57.operation_mode = "rom";
defparam ram_block1a57.port_a_address_clear = "none";
defparam ram_block1a57.port_a_address_width = 13;
defparam ram_block1a57.port_a_data_out_clear = "none";
defparam ram_block1a57.port_a_data_out_clock = "clock0";
defparam ram_block1a57.port_a_data_width = 1;
defparam ram_block1a57.port_a_first_address = 16384;
defparam ram_block1a57.port_a_first_bit_number = 9;
defparam ram_block1a57.port_a_last_address = 24575;
defparam ram_block1a57.port_a_logical_ram_depth = 65536;
defparam ram_block1a57.port_a_logical_ram_width = 24;
defparam ram_block1a57.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a57.ram_block_type = "auto";
defparam ram_block1a57.mem_init3 = "56AA552A954AAD56AA556AA556AA556AA554AAD55AAB556AAD55AAB554AAB554AAB554AAA555AAAD554AAA5556AAA5556AAAD555AAAA5554AAAA55552AAA95555AAAAB55554AAAAB55555AAAAAB555554AAAAAAD5555552AAAAAAA555555554AAAAAAAAAAD5555555555556AAAAAAAAAAAAAAAAAAAAAAAAAB555555555555555AAAAAAAAAAAAAAAAAAAAAAAAAA55555555555552AAAAAAAAA9555555552AAAAAAB5555554AAAAAA555555AAAAA955554AAAAB55556AAAAD5556AAAB5555AAAA5554AAA95552AAB5552AA9555AAAD556AA9556AA9556AA9552AAD55AAB556AA554AAD54AAD54AAD54AAD56AB552A954AA552A954AB55AA552AD56A956A956A956";
defparam ram_block1a57.mem_init2 = "A956AD52AD5AA54A956AD5AB54A952A54A952B56AD5A952A56AD4A95AB52B56A56A54AD4AD4AD4AD4AD4AD4A56A56A52B5295AD4AD6A5295AD4A52B5AD4A5295AD6B5AD6A5294A5294A52D6B5AD6B4A5294B5AD694A5AD294B5A52D694B5A52D694B4A5A52D29694B4B5A5A5AD2D2D2969696969696969696969696969696D2D2D2DA5A5B4B49696D2D25A4B49692D25B4B692D25B496D25B496D25B496DA4B6D25B692DB492DB4925B6924B6DA492DB692496DB6D24924B6DB6DB4924924924925B6DB6DB6DB6DB249249249249B6DB6D924924DB6D924936DB24936DB249B6C926DB24DB649B64936C936C93649B64DB24D926C9364DB26C9364D9364DB26C";
defparam ram_block1a57.mem_init1 = "9B26C9B264D9364D9B26C99364C9B364C9B364C99366CD9B366CD9B366CD9B3664C99B3664C99B3266CC99B33664CC99B336664CC9993336664CCC999933326666CCCCD9999933333366666664CCCCCCCCCC999999999999999999999999999999CCCCCCCCCCC6666666333333199998CCCCE66673331999CCCE666333999CCC66733199CCE6633198CC6633198CE673398CE67319CC67319CC67319CE6339CC67398C6739CC6319CE739CC6318C6318C6318C6318C739CE718C639CE718C738C639C639CE31CE31C639C638C718E71CE38C718E39C718E38C71C638E38C71C71C638E38E38E38E38E38E38E38E38E38E3C71C71C78E38E1C71E38E1C71E38F1";
defparam ram_block1a57.mem_init0 = "C78E1C70E3C70E3C78E1C38F1E3870E1C3870E1C3878F1E3C3870F1E1C3C7878F0F1E1E3C3C38787878F0F0F0F0F0F0F0F0F0F0F0F0F87878783C3C1E1E0F0F8783C3E1F0F8783C1F0F87C3E0F07C3E0F07C1F0F83E0F83E0F83E0F83E0F83E07C1F03E0FC1F03E07C0F81F03F07E07E0FC0FC0FC0FC0FC0FC0FC07E07F03F01F80FC07F01F80FE03F80FE03F807F01FE03FC07F807F00FF00FF007F807FC03FE00FF807FE00FF803FF003FE007FF003FF001FFC007FF001FFE001FFE001FFF0007FFE000FFFE0007FFF0000FFFF00007FFFE00003FFFFC00001FFFFF8000003FFFFFF80000000FFFFFFFFF800000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a81(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a81_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a81.clk0_core_clock_enable = "ena0";
defparam ram_block1a81.clk0_input_clock_enable = "ena0";
defparam ram_block1a81.clk0_output_clock_enable = "ena0";
defparam ram_block1a81.data_interleave_offset_in_bits = 1;
defparam ram_block1a81.data_interleave_width_in_bits = 1;
defparam ram_block1a81.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a81.init_file_layout = "port_a";
defparam ram_block1a81.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a81.operation_mode = "rom";
defparam ram_block1a81.port_a_address_clear = "none";
defparam ram_block1a81.port_a_address_width = 13;
defparam ram_block1a81.port_a_data_out_clear = "none";
defparam ram_block1a81.port_a_data_out_clock = "clock0";
defparam ram_block1a81.port_a_data_width = 1;
defparam ram_block1a81.port_a_first_address = 24576;
defparam ram_block1a81.port_a_first_bit_number = 9;
defparam ram_block1a81.port_a_last_address = 32767;
defparam ram_block1a81.port_a_logical_ram_depth = 65536;
defparam ram_block1a81.port_a_logical_ram_width = 24;
defparam ram_block1a81.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a81.ram_block_type = "auto";
defparam ram_block1a81.mem_init3 = "CC67319CC67319CC67319CC67319CC67319CC67319CC673198CE63398CE63398CE63398CE63398CE67319CC67319CC67319CC673398CE63398CE63399CC67319CC673198CE63398CE63319CC67319CCE63398CE67319CC673398CE63319CC673398CE63319CC663398CE67319CCE63399CC673398CC673198CE67319CCE63319CCE63319CCE63319CCE63319CCE63319CCE673198CC673398CC663399CCE673198CC663399CCE673398CC6633198CC6633198CC6633198CC6633198CC6633198CC6673399CCE6733198CC6673399CCC6633399CCC6633399CCC66333998CC66733199CCE66333998CCE66333998CCE66333199CCC667333998CCE667331998CC";
defparam ram_block1a81.mem_init2 = "C667333999CCCE667333999CCCE6673331998CCC66673331998CCCE66633339998CCCC666733339998CCCC6666333319999CCCCE66663333399998CCCCC6666633333199999CCCCCC6666673333339999998CCCCCCC666666633333333199999999CCCCCCCCCC6666666666673333333333333319999999999999999999999CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC9999999999999999999999B3333333333333266666666664CCCCCCCCD99999999B33333326666664CCCCCC999999333332666664CCCCD9999B333366666CCCC9999B33326666CCCD999B3336666CCCD9993332666CCC999B332666CCD999332666CCD99B33666CCD99B33666CC9";
defparam ram_block1a81.mem_init1 = "9933666CC99933664CC99B3266CC99B3266CC99B3664CD993266CD993266CD993266CD9B3664C993266CD9B366CD9B366CD9B366CD93264C99366CD9B264C9B366C99366C99366C99366C99364C9B264D9326C99364D9B26C9B364D9364D9326C9B26C9B26C9B26C9B26C9B26D9364D93649B26C9B64D926C9B24D926C9B64DB26D936C9B64DB24D926D926C936C936C936C936C936C936C926D926DB24DB649B6C926DB249B6C926DB24936D9249B6D9249B6D924936DB64924DB6DB249249B6DB6D924924936DB6DB6DB24924924924924924924924924924924924924924924B6DB6DB6DB4924924B6DB6DA492496DB6D24925B6DA4925B6D2492DB6924B6";
defparam ram_block1a81.mem_init0 = "D2496DA492DB492DB492DB492DB496DA496D24B692DB496D25B692DA4B692DA4B692D25B496D2DA4B696D2DA4B49692D25A4B49692D2DA5B4B4969692D2DA5A5A4B4B4B696969696D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D29696969694B4B4B5A5A52D2D29694B4B5A5AD2D696B4A5A52D694B5A5AD296B5A52D694A5AD294B5AD294B5AD694A5296B5AD6B4A5294A5294A5294A5294A5294A56B5AD6B5294A56B5A94A56B5A94AD6A52B5A94AD6A56B52B5A95A94AD4AD4AD4A56A56A56A56AD4AD4AD4A95A952B52A56A54AD5AB52A56AD5A952A54A952A54A952A54A952A55AB56A952AD5AA54AB54A956A956A956A956A954AB54AA55AAD52A954AB55AAD";

cyclonev_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "rom";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "clock0";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 8191;
defparam ram_block1a9.port_a_logical_ram_depth = 65536;
defparam ram_block1a9.port_a_logical_ram_width = 24;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init3 = "6AB55AA552A956AB54AA55AA552AD52AD52AD52AD52A55AA54AB56A952AD5AB54A952A54A952A54A952A54A952B56AD4A95AB56A54AD4A95A952B52A56A56A56AD4AD4AD4AD4A56A56A56A52B52B5A95AD4AD6A52B5A94AD6A52B5AD4A52B5AD4A5295AD6B5AD4A5294A5294A5294A5294A5294A5AD6B5AD294A52D6B5A5296B5A5296B4A52D694B5AD296B4B5A52D694B4A5AD2D696B4B5A5A52D2969694B4B5A5A5A52D2D2D2D296969696969696969696969696969696D2D2D2D2DA5A5A4B4B4B69692D2D25A5B4B69692D25A4B49692D25A4B696D2DA4B696D25B49692DA4B692DA4B692DB496D25B692DA496D24B6D25B6925B6925B6925B6924B6D2496";
defparam ram_block1a9.mem_init2 = "DA492DB692496DB4924B6DB492496DB6D24924B6DB6DA4924925B6DB6DB6DA49249249249249249249249249249249249249249249B6DB6DB6D924924936DB6DB249249B6DB64924DB6D924936DB24936DB24936D9249B6C926DB249B6C926DB24DB649B6C936C926D926D926D926D926D926D926C936C93649B64DB26D936C9B64DB26C93649B26C9364DB26C9B24D9364D936C9B26C9B26C9B26C9B26C9B26C99364D9364D9B26C9B364D9326C99364C9B264D9326CD9326CD9326CD9326CD9B264C9B366CD93264C99366CD9B366CD9B366CD9B366CC993264CD9B366CC993366CC993366CC9933664CD9B3266CC99B3266CC99B32664CD9933266CCD9933";
defparam ram_block1a9.mem_init1 = "266CCD99B33666CCD99B33666CCC999333666CCC999B332666CCC99993336666CCCD999B3336666CCCC9999B33326666CCCCD9999B3333666664CCCCC9999993333326666664CCCCCC9999999B333333336666666664CCCCCCCCCC99999999999999B33333333333333333333326666666666666666666666666666666666666673333333333333333333333199999999999999CCCCCCCCCCCC666666666733333333199999998CCCCCCC66666663333333999999CCCCCC66666733333199998CCCCC666663333399998CCCCE6667333319998CCCC666633339999CCCC666633339998CCCE6663331999CCCC6663331999CCCE667333999CCCE667333999CCC6";
defparam ram_block1a9.mem_init0 = "66333199CCCE66333999CCC667331998CCE66333998CCE66333998CCE6733199CCC66333998CC66733998CC66733998CC6673399CCC6633199CCE673399CCC6633198CC6633198CC6633198CC6633198CC6633198CC663399CCE673398CC663319CCE673398CC663399CC663319CCE673198CE673198CE673198CE673198CE673198CE67319CCE63319CC663399CC673398CE67319CCE63398CC673198CE63399CC673198CE63399CC67319CCE63398CE67319CC673198CE63398CE63319CC67319CC673398CE63398CE63399CC67319CC67319CC67319CCE63398CE63398CE63398CE63398CE63319CC67319CC67319CC67319CC67319CC67319CC67319CC66";

cyclonev_ram_block ram_block1a33(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a33_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a33.clk0_core_clock_enable = "ena0";
defparam ram_block1a33.clk0_input_clock_enable = "ena0";
defparam ram_block1a33.clk0_output_clock_enable = "ena0";
defparam ram_block1a33.data_interleave_offset_in_bits = 1;
defparam ram_block1a33.data_interleave_width_in_bits = 1;
defparam ram_block1a33.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a33.init_file_layout = "port_a";
defparam ram_block1a33.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a33.operation_mode = "rom";
defparam ram_block1a33.port_a_address_clear = "none";
defparam ram_block1a33.port_a_address_width = 13;
defparam ram_block1a33.port_a_data_out_clear = "none";
defparam ram_block1a33.port_a_data_out_clock = "clock0";
defparam ram_block1a33.port_a_data_width = 1;
defparam ram_block1a33.port_a_first_address = 8192;
defparam ram_block1a33.port_a_first_bit_number = 9;
defparam ram_block1a33.port_a_last_address = 16383;
defparam ram_block1a33.port_a_logical_ram_depth = 65536;
defparam ram_block1a33.port_a_logical_ram_width = 24;
defparam ram_block1a33.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.ram_block_type = "auto";
defparam ram_block1a33.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000003FFFFFFFFE00000003FFFFFF8000003FFFFF000007FFFF80000FFFFC0001FFFE0001FFFC000FFFE000FFFC001FFF000FFF000FFF001FFC007FF001FF801FFC00FF801FF803FE00FFC03FE00FF807FC03FC01FE01FE01FC03FC07F80FF01FC03F80FE03F80FE03F01FC07E03F01F81FC0FC07E07E07E07E07E07E07E0FC0FC1F81F03E07C0F81F07E0F81F07C0F83E0F83E0F83E0F83E0F83E1F07C1E0F87C1E0F87C3E1F0783C3E1F0F8783C3E1E0F0F078783C3C3C3E1E1E1E1E1E1E1E1E1E1E1E1E3C3C3C387878F0F1E1E3C3C7870F1E1C3878F1E3C3870E1C3870E1C38F1E3870E3C78E1C78E1C70E3C7";
defparam ram_block1a33.mem_init2 = "1E38F1C70E38F1C70E38E3C71C71C78E38E38E38E38E38E38E38E38E38E38C71C71C638E38C71C638E31C738E31C638E71CE31C638C738C718E718E738C738C639C631CE738C631CE739C6318C6318C6318C6318C6739CE7318C6739CC6339CC67398CE7319CC67319CC67319CCE63399CCE633198CC6633198CCE6733199CCC667333998CCCE6673331999CCCCE6666333331999998CCCCCCC6666666666733333333333333333333333333333266666666664CCCCCCD9999993333366666CCCC999933326664CCD999332664CCD99B32664CD99B3266CC99B3264CD9B3264CD9B366CD9B366CD9B366CD93264D9B264D9B264D9326C9B364D9364C9B26C9B2";
defparam ram_block1a33.mem_init1 = "6C9B64D9364D926C9B64D926C93649B64DB24D926D926D924DB24DB649B6C926DB249B6D9249B6D924936DB64924936DB6DB249249249249B6DB6DB6DB6DB4924924924925B6DB6DA492496DB6D2492DB6924B6DA492DB4925B6925B692DB496DA4B6D25B496D25B496D25B49692DA5B49692D25A4B49696D2D25A5B4B4B6969696D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2969696B4B4B5A5A52D29694B4A5A52D694B5A52D694B5A5296B4A52D6B5A5294A5AD6B5AD694A5294A5294AD6B5AD6B5294A56B5A94A56B5294AD6A56B5295A94AD4AD4A56A56A56A56A56A56A54AD4AD5A95AB52A56AD4A952B56AD5A952A54A952A55AB56AD52A54AB56A956AD52A";
defparam ram_block1a33.mem_init0 = "D52AD52AD52AD56A954AB55AA552A954AA552A955AAD56AA556AA556AA556AA554AAD55AAB556AA9552AAD552AAD552AAD556AAB5552AA9555AAA95552AAA5554AAAB5555AAAAD5556AAAAD5555AAAAA555552AAAAB555554AAAAAA5555555AAAAAAA9555555552AAAAAAAAA95555555555554AAAAAAAAAAAAAAAAAAAAAAAAAB555555555555555AAAAAAAAAAAAAAAAAAAAAAAAAAD5555555555556AAAAAAAAAA555555554AAAAAAA95555556AAAAAA555555AAAAAB55555AAAAA55555AAAAB55552AAA95554AAAA5554AAAB5556AAAD554AAAD554AAA5556AAB554AAA555AAA555AAA555AAB556AAD55AAB556AA554AAD54AAD54AAD54AAD56AA552A954AAD5";

cyclonev_ram_block ram_block1a106(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a106_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a106.clk0_core_clock_enable = "ena0";
defparam ram_block1a106.clk0_input_clock_enable = "ena0";
defparam ram_block1a106.clk0_output_clock_enable = "ena0";
defparam ram_block1a106.data_interleave_offset_in_bits = 1;
defparam ram_block1a106.data_interleave_width_in_bits = 1;
defparam ram_block1a106.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a106.init_file_layout = "port_a";
defparam ram_block1a106.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a106.operation_mode = "rom";
defparam ram_block1a106.port_a_address_clear = "none";
defparam ram_block1a106.port_a_address_width = 13;
defparam ram_block1a106.port_a_data_out_clear = "none";
defparam ram_block1a106.port_a_data_out_clock = "clock0";
defparam ram_block1a106.port_a_data_width = 1;
defparam ram_block1a106.port_a_first_address = 32768;
defparam ram_block1a106.port_a_first_bit_number = 10;
defparam ram_block1a106.port_a_last_address = 40959;
defparam ram_block1a106.port_a_logical_ram_depth = 65536;
defparam ram_block1a106.port_a_logical_ram_width = 24;
defparam ram_block1a106.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a106.ram_block_type = "auto";
defparam ram_block1a106.mem_init3 = "B3266CC99B3264CD993366CC99B3664C99B3664C99B366CC993264CD9B366CD993264C993264C993264C993264D9B366CD93264C99366CD93264D9B364C9B364C99366C99366C9B364C9B364D9B26CD9366C9B364D9326C9B364D9366C9B26C99364D9364D9366C9B26C9B26C9B26C9B26C9B26C9364D9364D93649B26C9B24D9364DB26C9B64D926C9B24D926C9B64D926C93649B24D926C93649B24DB26D926C936C9B649B649B24DB24DB24DB24DB24DB24DB24DB24DB649B649B6C936C926D924DB249B64936D924DB249B6C926DB249B6C924DB64936DB249B6D924DB6C924DB6C924DB6D9249B6DB24936DB649249B6DB24924DB6DB24924DB6DB64924";
defparam ram_block1a106.mem_init2 = "936DB6DB24924926DB6DB6D9249249249B6DB6DB6DB6C924924924924924936DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6D24924924924924925B6DB6DB6DB6D2492492496DB6DB6DA4924925B6DB6DA492492DB6DB492492DB6DB492496DB6D24925B6DB4924B6DB4924B6DB4924B6DB4925B6DA492DB6924B6DA492DB6924B6DA492DB4925B6924B6D2496DA496DA492DB492DB492DB492DB492DB492DA496DA496D24B6D25B6925B492DA496D24B6925B496DA4B6925B496DA4B692DB496D25B496DA4B692DA4B692DA4B692DA4B692DA4B692DA4B696D25B496D25A4B692DA5B496D25A4B696D25B4B692D25B4B692D25B4B696D25A4B49692DA5";
defparam ram_block1a106.mem_init1 = "B4B696D2DA5B4B696D2DA5B4B696D2DA5A4B49692D2DA5B4B49692D2DA5A4B4B69692D2DA5A4B4B69692D2D25A5B4B4B69696D2D2DA5A5B4B4B6969692D2D2DA5A5A4B4B4B496969692D2D2D2DA5A5A5A5B4B4B4B4B69696969696D2D2D2D2D2D2D2DA5A5A5A5A5A5A5A5A5A5A4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4A5A5A5A5A5A5A5A5A5A5A5A52D2D2D2D2D2D2D6969696969694B4B4B4B4A5A5A5A5A52D2D2D2D6969696B4B4B4B5A5A5A52D2D2D6969694B4B4A5A5A5AD2D2D69696B4B4B5A5A52D2D29696B4B4A5A5A52D2D69694B4B5A5AD2D29696B4B4A5A52D2D696B4B4A5A52D29696B4B5A5AD2D696B4B5A5AD2D696B4B5A5AD2D696B";
defparam ram_block1a106.mem_init0 = "4B5A52D29694B4A5AD2D696B4A5A52D296B4B5A52D296B4B5A52D296B4A5A52D696B4A5AD2D694B5A52D296B4A5AD2D694B5A52D696B4A5AD296B4A5AD29694B5A52D694B5A52D694B5A52D694B5A52D694B5A52D694B5AD296B4A5AD296B4A5AD694B5A52D694B5AD296B4A5AD694B5A52D6B4A5AD294B5A52D6B4A5AD294B5A52D6B4A5AD694B5A5296B4A52D694A5AD294B5A5296B4A52D694A5AD294B5AD296B5A52D6B4A52D694A5AD694B5AD294B5A5296B5A52D6B4A52D6B4A5AD694A5AD694A5AD294B5AD294B5AD296B5A5296B5A5296B5A5296B4A52D6B4A52D6B4A52D6B4A52D6B4A5AD694A5AD694A5AD694A5AD694A5AD694A5AD694A5AD694A";

cyclonev_ram_block ram_block1a130(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a130_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a130.clk0_core_clock_enable = "ena0";
defparam ram_block1a130.clk0_input_clock_enable = "ena0";
defparam ram_block1a130.clk0_output_clock_enable = "ena0";
defparam ram_block1a130.data_interleave_offset_in_bits = 1;
defparam ram_block1a130.data_interleave_width_in_bits = 1;
defparam ram_block1a130.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a130.init_file_layout = "port_a";
defparam ram_block1a130.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a130.operation_mode = "rom";
defparam ram_block1a130.port_a_address_clear = "none";
defparam ram_block1a130.port_a_address_width = 13;
defparam ram_block1a130.port_a_data_out_clear = "none";
defparam ram_block1a130.port_a_data_out_clock = "clock0";
defparam ram_block1a130.port_a_data_width = 1;
defparam ram_block1a130.port_a_first_address = 40960;
defparam ram_block1a130.port_a_first_bit_number = 10;
defparam ram_block1a130.port_a_last_address = 49151;
defparam ram_block1a130.port_a_logical_ram_depth = 65536;
defparam ram_block1a130.port_a_logical_ram_width = 24;
defparam ram_block1a130.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a130.ram_block_type = "auto";
defparam ram_block1a130.mem_init3 = "00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFC0000000000003FFFFFFFFFF8000000000FFFFFFFFE00000001FFFFFFF0000000FFFFFFE000000FFFFFF000001FFFFF800001FFFFE00000FFFFE00003FFFF00003FFFF00007FFFC0001FFFE0001FFFC0007FFF0001FFFC000FFFC000FFFC001FFF8003FFE001FFF0007FF8007FF8007FF8007FF000FFE001FFC007FF001FF800FFE007FF003FF003FF003FF003FF003FE007FE00FF801FF007FC01FF803FC01FF007FC03FE00FF007F803FC03FC01FE01FE01FE01FE01FE01FE03FC03FC07F80FF01FE03FC07F80FE01FC07F01FC03F80FE03F80FE07F01FC07F03F80FE07F01F80FC07";
defparam ram_block1a130.mem_init2 = "E03F01F80FC0FE07F03F03F81F81F80FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0F81F81F83F03F07E07C0FC1F83F03E07C0F81F03E07C0F83F07C0F81F07C0F83F07C1F83E0F83F07C1F07C1F83E0F83E0F83E0F83E0F87C1F07C1F0783E0F83C1F0783E0F07C1E0F87C1E0F87C1E0F07C3E1F0F83C1E0F0783C1E0F0F87C3E1E0F0787C3C1E1F0F0787C3C1E1E0F0F078783C3C3E1E1E1F0F0F0F078787878787C3C3C3C3C3C3C3C3C3C3C3C3C3C3C387878787878F0F0F0E1E1E1E3C3C387878F0F0E1E1C3C387870F1E1E3C3878F0E1E3C3878F1E1C3C78F0E1C3C78F1E3C3870E1C3870E1C3870E1C3870E1C3871E3C78E1C3871E3C70E3C78E1C78F1C38F1C3";
defparam ram_block1a130.mem_init1 = "8F1C78E1C78E1C70E3871E38F1C78E3871C38E3C71E38E1C71C38E3871C70E38E3C71C71E38E38E1C71C71C78E38E38E38E3C71C71C71C71C71C71C71C71C71C71C71C71C638E38E38E38E71C71C71CE38E38C71C71CE38E39C71C638E31C718E38C71C638E71C638E71C638E71CE39C718E31C638C718E71CE39C638C738E718E71CE31CE31CE31CE31CE31CE31CE31CE718E738C739C639CE318E738C639CE718C639CE718C639CE738C6318C639CE739CE739CE718C6318C6318CE739CE739CE7398C6318C6739CE7318C6739CE6318CE7318C67398C67398C67398C67318CE6319CC63398CE7319CC67319CE63398CE63399CC67319CC673398CE67319CC";
defparam ram_block1a130.mem_init0 = "E63319CCE633198CE673399CC6633198CC6633199CCE6733998CC66733998CC66733199CCC66733199CCCE66333199CCCE667333999CCCE6663331999CCCC666733339999CCCCE6667333319999CCCCC66666333333999998CCCCCC66666663333333199999999CCCCCCCCCCE6666666666667333333333333333333333333339999999999999993333333333333333333333333366666666666664CCCCCCCCCC999999999333333326666664CCCCCC99999933333266666CCCCC999993333266664CCCD999933336666CCCD999B3336666CCC99993336664CCD999333666CCC999333666CCD99B33666CCD99B33666CC99933666CC99933664CC99B3266CC99";

cyclonev_ram_block ram_block1a154(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a154_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a154.clk0_core_clock_enable = "ena0";
defparam ram_block1a154.clk0_input_clock_enable = "ena0";
defparam ram_block1a154.clk0_output_clock_enable = "ena0";
defparam ram_block1a154.data_interleave_offset_in_bits = 1;
defparam ram_block1a154.data_interleave_width_in_bits = 1;
defparam ram_block1a154.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a154.init_file_layout = "port_a";
defparam ram_block1a154.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a154.operation_mode = "rom";
defparam ram_block1a154.port_a_address_clear = "none";
defparam ram_block1a154.port_a_address_width = 13;
defparam ram_block1a154.port_a_data_out_clear = "none";
defparam ram_block1a154.port_a_data_out_clock = "clock0";
defparam ram_block1a154.port_a_data_width = 1;
defparam ram_block1a154.port_a_first_address = 49152;
defparam ram_block1a154.port_a_first_bit_number = 10;
defparam ram_block1a154.port_a_last_address = 57343;
defparam ram_block1a154.port_a_logical_ram_depth = 65536;
defparam ram_block1a154.port_a_logical_ram_width = 24;
defparam ram_block1a154.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a154.ram_block_type = "auto";
defparam ram_block1a154.mem_init3 = "3266CC99B32664CD9933266CCD9933266CCD99B33666CCD99B33666CCD999332666CCD9993336664CCD9993332666CCCD999B3336666CCCD9999333366664CCCC999993333266666CCCCC9999993333326666664CCCCCC9999999933333333266666666664CCCCCCCCCCCCD9999999999999999999999999933333333333333399999999999999999999999999CCCCCCCCCCCCCE66666666673333333319999998CCCCCCC666666333333999998CCCCC66667333319999CCCCE666733339999CCCC66673331998CCCE667333999CCCE667331998CCE66733199CCC66733199CCC6633399CCC6633399CCE6733198CC6633198CC673399CCE633198CE673198CE";
defparam ram_block1a154.mem_init2 = "67319CCE63399CC67319CC673398CE63398CE7319CC67319CE63398C67318CE6319CC6339CC6339CC6339CC6319CE6318CE739CC6319CE739CC6318C6339CE739CE739CE6318C6318C631CE739CE739CE738C6318C639CE738C631CE738C631CE738C639CE318E738C739C639CE31CE718E718E718E718E718E718E718E71CE31CE39C638C738E71CE31C638C718E31C738E71CE38C71CE38C71CE38C71C638E31C718E38C71C738E38E71C71C638E38E71C71C71CE38E38E38E38C71C71C71C71C71C71C71C71C71C71C71C71C78E38E38E38E3C71C71C70E38E38F1C71C78E38E1C71C38E3871C70E38F1C78E3871C38E3C71E38F1C38E1C70E3C70E3C71E3";
defparam ram_block1a154.mem_init1 = "871E3871E3C70E3C78E1C78F1C3870E3C78F1C3870E1C3870E1C3870E1C3870E1C3878F1E3C7870E1E3C7870F1E3C3878F0E1E3C3878F0F1E1C3C387870F0E1E1E3C3C387878F0F0F0E1E1E1E3C3C3C3C3C3878787878787878787878787878787C3C3C3C3C3C1E1E1E1F0F0F0F878783C3C1E1E0F0F0787C3C1E1F0F0787C3C1E0F0F87C3E1E0F0783C1E0F0783E1F0F87C1E0F07C3E0F07C3E0F07C1E0F83C1F0783E0F83C1F07C1F07C3E0F83E0F83E0F83E0F83F07C1F07C1F83E0F83F07C1F83E07C1F03E07C1F83E07C0F81F03E07C0F81F83F07E07C0FC1F81F83F03F03E07E07E07E07E07E07E07E07E07E07E03F03F03F81F81FC0FE07E03F01F80F";
defparam ram_block1a154.mem_init0 = "C07E03F01FC0FE03F81FC07F01FC0FE03F80FE03F807F01FC07F00FE03FC07F80FF01FE03FC07F807F80FF00FF00FF00FF00FF00FF007F807F803FC01FE00FF807FC01FF007F803FF007FC01FF003FE00FFC00FF801FF801FF801FF801FF801FFC00FFE003FF001FFC007FF000FFE001FFC003FFC003FFC003FFC001FFF000FFF8003FFF0007FFE0007FFE0007FFF0001FFFC0007FFF0000FFFF00007FFFC0001FFFF80001FFFF80000FFFFE00000FFFFF000003FFFFF000001FFFFFE000000FFFFFFE0000001FFFFFFF00000000FFFFFFFFE0000000003FFFFFFFFFF80000000000007FFFFFFFFFFFFFFFF80000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a178(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a178_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a178.clk0_core_clock_enable = "ena0";
defparam ram_block1a178.clk0_input_clock_enable = "ena0";
defparam ram_block1a178.clk0_output_clock_enable = "ena0";
defparam ram_block1a178.data_interleave_offset_in_bits = 1;
defparam ram_block1a178.data_interleave_width_in_bits = 1;
defparam ram_block1a178.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a178.init_file_layout = "port_a";
defparam ram_block1a178.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a178.operation_mode = "rom";
defparam ram_block1a178.port_a_address_clear = "none";
defparam ram_block1a178.port_a_address_width = 13;
defparam ram_block1a178.port_a_data_out_clear = "none";
defparam ram_block1a178.port_a_data_out_clock = "clock0";
defparam ram_block1a178.port_a_data_width = 1;
defparam ram_block1a178.port_a_first_address = 57344;
defparam ram_block1a178.port_a_first_bit_number = 10;
defparam ram_block1a178.port_a_last_address = 65535;
defparam ram_block1a178.port_a_logical_ram_depth = 65536;
defparam ram_block1a178.port_a_logical_ram_width = 24;
defparam ram_block1a178.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a178.ram_block_type = "auto";
defparam ram_block1a178.mem_init3 = "A52D6B4A52D6B4A52D6B4A52D6B4A52D6B4A52D6B4A52D6B4A5AD694A5AD694A5AD694A5AD694A5AD294B5AD294B5AD294B5AD296B5A5296B5A5296B4A52D6B4A52D6B4A5AD694A5AD694B5AD294B5A5296B5A52D6B4A52D694A5AD694B5AD296B5A5296B4A52D694A5AD294B5A5296B4A52D694A5AD294B5A52D6B4A5AD694B5A5296B4A5AD694B5A5296B4A5AD694B5A52D6B4A5AD296B5A52D694B5A52D6B4A5AD296B4A5AD296B5A52D694B5A52D694B5A52D694B5A52D694B5A52D694B5A52D296B4A5AD296B4A5AD2D694B5A52D696B4A5AD29694B5A52D696B4A5AD2D694B4A5AD29694B5A5AD29694B5A5AD29694B4A5AD2D696B4A5A52D29694B5A5";
defparam ram_block1a178.mem_init2 = "AD2D696B4B5A5AD2D696B4B5A5AD2D696B4B5A5AD2D29694B4A5A5AD2D69694B4A5A5AD2D29696B4B5A5A52D2D69694B4B4A5A5AD2D2969694B4B5A5A5AD2D2D69696B4B4B4A5A5A52D2D2D6969694B4B4B5A5A5A5AD2D2D2D696969694B4B4B4B4A5A5A5A5A52D2D2D2D2D2D696969696969694B4B4B4B4B4B4B4B4B4B4B4A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A4B4B4B4B4B4B4B4B4B4B4B696969696969696D2D2D2D2D2DA5A5A5A5B4B4B4B4B696969692D2D2D25A5A5A4B4B4B6969692D2D2DA5A5B4B4B69696D2D2DA5A5B4B4969692D2DA5A4B4B69692D2DA5A4B4B69692D25A5B4B69692D25A4B4B696D2DA5B4B696D2DA5B4B696D2DA5B";
defparam ram_block1a178.mem_init1 = "4B692D25A4B496D2DA5B49692DA5B49692DA5B496D2DA4B496D25B4B692DA4B496D25B496D2DA4B692DA4B692DA4B692DA4B692DA4B692DA4B6D25B496D25B692DA4B6D25B492DA4B6D25B492DA496D24B6925B492DB496DA496D24B6D24B6925B6925B6925B6925B6925B6924B6D24B6D2496DA492DB4925B6924B6DA492DB6924B6DA492DB6924B6DB4925B6DA4925B6DA4925B6DA4925B6DB492496DB6D24925B6DB6924925B6DB6924924B6DB6DB4924924B6DB6DB6D2492492496DB6DB6DB6DB492492492492492496DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6D924924924924924926DB6DB6DB6DB24924924936DB6DB6C9249249B6DB6D92";
defparam ram_block1a178.mem_init0 = "4924DB6DB649249B6DB649249B6DB24924DB6D9249B6DB24936DB64926DB64926DB64936DB249B6D924DB64926DB249B6C926DB249B64936D924DB249B64936C926D926DB24DB24DB649B649B649B649B649B649B649B649B24DB24DB26D926C936C9B649B24D926C93649B24D926C9364DB26C93649B26C9364DB26C9B64D93649B26C9B24D9364D9364D926C9B26C9B26C9B26C9B26C9B26CD9364D9364D9326C9B26CD9364D9B26C99364D9B26CD9366C9B364D9B264D9B26CD9326CD93264D9B264D9B364C99366CD93264C99366CD9B364C993264C993264C993264C993366CD9B3664C993266CD9B3264CD9B3264CD9B3266CD9933664C99B3266CC99B";

cyclonev_ram_block ram_block1a58(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a58_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a58.clk0_core_clock_enable = "ena0";
defparam ram_block1a58.clk0_input_clock_enable = "ena0";
defparam ram_block1a58.clk0_output_clock_enable = "ena0";
defparam ram_block1a58.data_interleave_offset_in_bits = 1;
defparam ram_block1a58.data_interleave_width_in_bits = 1;
defparam ram_block1a58.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a58.init_file_layout = "port_a";
defparam ram_block1a58.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a58.operation_mode = "rom";
defparam ram_block1a58.port_a_address_clear = "none";
defparam ram_block1a58.port_a_address_width = 13;
defparam ram_block1a58.port_a_data_out_clear = "none";
defparam ram_block1a58.port_a_data_out_clock = "clock0";
defparam ram_block1a58.port_a_data_width = 1;
defparam ram_block1a58.port_a_first_address = 16384;
defparam ram_block1a58.port_a_first_bit_number = 10;
defparam ram_block1a58.port_a_last_address = 24575;
defparam ram_block1a58.port_a_logical_ram_depth = 65536;
defparam ram_block1a58.port_a_logical_ram_width = 24;
defparam ram_block1a58.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a58.ram_block_type = "auto";
defparam ram_block1a58.mem_init3 = "CD9933664CD99B3266CCD9933266CCD99332664CC999332664CC999332666CCD999332666CCC999B332666CCCD99933326664CCC999933326666CCCC9999B333366666CCCCD9999933333666666CCCCCD999999B33333366666666CCCCCCCCD9999999999B333333333333266666666666666666666666666CCCCCCCCCCCCCCC66666666666666666666666666333333333333319999999998CCCCCCCCE66666673333333999999CCCCCC6666673333399998CCCCE6666333319998CCCC666633339998CCCE6673331998CCC6663331998CCE667331998CCE66333998CCE6633399CCC6633399CCC6633198CCE673399CCE673398CC663319CCE673198CE6731";
defparam ram_block1a58.mem_init2 = "98CE63319CC663398CE63398CC67319CC67318CE63398CE6319CC67398CE7319CE6339CC6339CC6339CC6339CE6319CE7318C6339CE6318C6339CE739CC6318C6318C6319CE739CE739CE318C6318C6318C739CE739C6318C739CE318C739CE318C739C631CE718C738C639C631CE318E718E718E718E718E718E718E718E31CE31C639C738C718E31CE39C738E71CE38C718E31C738E31C738E31C738E39C71CE38E71C738E38C71C718E38E39C71C718E38E38E31C71C71C71C738E38E38E38E38E38E38E38E38E38E38E38E3871C71C71C71C38E38E38F1C71C70E38E3871C71E38E3C71C78E38F1C70E38F1C78E3C71C38E1C70E3C71E38F1C38F1C38E1C";
defparam ram_block1a58.mem_init1 = "78E1C78E1C38F1C3871E3870E3C78F1C3870E3C78F1E3C78F1E3C78F1E3C78F1E3C7870E1C3878F1E1C3878F0E1C3C7870F1E1C3C7870F0E1E3C3C7878F0F1E1E1C3C3C787870F0F0F1E1E1E1C3C3C3C3C3C7878787878787878787878787878783C3C3C3C3C3E1E1E1E0F0F0F078787C3C3E1E1F0F0F8783C3E1E1F0F8783C3E1F0F0783C1E1F0F87C3E1F0F87C1E0F0783E1F0F83C1F0F83C1F0F83E1F07C3E0F87C1F07C3E0F83E0F83C1F07C1F07C1F07C1F07C0F83E0F83E07C1F07C0F83E07C1F83E0FC1F03E07C1F83F07E0FC1F83F07E07C0F81F83F03E07E07C0FC0FC1F81F81F81F81F81F81F81F81F81F81FC0FC0FC07E07E03F01F81FC0FE07F0";
defparam ram_block1a58.mem_init0 = "3F81FC0FE03F01FC07E03F80FE07F01FC07F01FC07F80FE03F80FF01FC03F807F00FE01FC03F807F807F00FF00FF00FF00FF00FF00FF807F807FC03FE01FF007F803FE00FF807FC00FF803FE00FFC01FF003FF007FE007FE007FE007FE007FE003FF001FFC00FFE003FF800FFF001FFE003FFC003FFC003FFC003FFE000FFF0007FFC000FFF8001FFF8001FFF8000FFFE0003FFF8000FFFF0000FFFF80003FFFE00007FFFE00007FFFF00001FFFFF00000FFFFFC00000FFFFFE000001FFFFFF0000001FFFFFFE0000000FFFFFFFF000000001FFFFFFFFFC00000000007FFFFFFFFFFFF800000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a82(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a82_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a82.clk0_core_clock_enable = "ena0";
defparam ram_block1a82.clk0_input_clock_enable = "ena0";
defparam ram_block1a82.clk0_output_clock_enable = "ena0";
defparam ram_block1a82.data_interleave_offset_in_bits = 1;
defparam ram_block1a82.data_interleave_width_in_bits = 1;
defparam ram_block1a82.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a82.init_file_layout = "port_a";
defparam ram_block1a82.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a82.operation_mode = "rom";
defparam ram_block1a82.port_a_address_clear = "none";
defparam ram_block1a82.port_a_address_width = 13;
defparam ram_block1a82.port_a_data_out_clear = "none";
defparam ram_block1a82.port_a_data_out_clock = "clock0";
defparam ram_block1a82.port_a_data_width = 1;
defparam ram_block1a82.port_a_first_address = 24576;
defparam ram_block1a82.port_a_first_bit_number = 10;
defparam ram_block1a82.port_a_last_address = 32767;
defparam ram_block1a82.port_a_logical_ram_depth = 65536;
defparam ram_block1a82.port_a_logical_ram_width = 24;
defparam ram_block1a82.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a82.ram_block_type = "auto";
defparam ram_block1a82.mem_init3 = "5AD294B5AD294B5AD294B5AD294B5AD294B5AD294B5AD294B5A5296B5A5296B5A5296B5A5296B5A52D6B4A52D6B4A52D6B4A52D694A5AD694A5AD694B5AD294B5AD294B5A5296B5A5296B4A52D6B4A5AD694A5AD294B5AD296B5A5296B4A52D694A5AD694B5AD296B5A52D6B4A5AD694B5AD296B5A52D6B4A5AD294B5A5296B4A5AD694B5A5296B4A5AD694B5A5296B4A5AD294B5A52D694A5AD296B4A5AD294B5A52D694B5A52D694A5AD296B4A5AD296B4A5AD296B4A5AD296B4A5AD296B4A5AD2D694B5A52D694B5A52D296B4A5AD29694B5A52D696B4A5AD29694B5A52D296B4B5A52D696B4A5A52D696B4A5A52D696B4B5A52D29694B5A5AD2D694B4A5A";
defparam ram_block1a82.mem_init2 = "52D29694B4A5A52D29694B4A5A52D29694B4A5A52D2D696B4B5A5A52D29696B4B5A5A52D2D69694B4A5A5AD2D29696B4B4B5A5A52D2D69696B4B4A5A5A52D2D2969694B4B4B5A5A5AD2D2D2969696B4B4B4A5A5A5A52D2D2D296969696B4B4B4B4B5A5A5A5A5AD2D2D2D2D2D296969696969696B4B4B4B4B4B4B4B4B4B4B4B5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5B4B4B4B4B4B4B4B4B4B4B49696969696969692D2D2D2D2D25A5A5A5A4B4B4B4B496969696D2D2D2DA5A5A5B4B4B4969696D2D2D25A5A4B4B4969692D2D25A5A4B4B69696D2D25A5B4B49696D2D25A5B4B49696D2DA5A4B49696D2DA5B4B49692D25A4B49692D25A4B49692D25A4";
defparam ram_block1a82.mem_init1 = "B496D2DA5B4B692D25A4B696D25A4B696D25A4B692D25B4B692DA4B496D25B4B692DA4B692D25B496D25B496D25B496D25B496D25B496D25B492DA4B692DA496D25B492DA4B6D25B492DA4B6D25B692DB496DA4B6D24B6925B692DB492DB496DA496DA496DA496DA496DA496DB492DB492DB6925B6D24B6DA496DB4925B6D2496DB4925B6D2496DB4924B6DA4925B6DA4925B6DA4925B6DA4924B6DB692492DB6DA492496DB6DA492496DB6DB4924924B6DB6DB492492492DB6DB6DB6924924924924B6DB6DB6DB6DB6DB6924924924924924924924924924924924924924924926DB6DB6DB6DB6DB6D924924924924DB6DB6DB6C924924936DB6DB64924926D";
defparam ram_block1a82.mem_init0 = "B6DB249249B6DB649249B6DB64924DB6DB24926DB64924DB6C9249B6D9249B6D9249B6C924DB64926DB249B6D924DB64936D924DB649B6C926DB24DB649B6C936D926D924DB24DB249B649B649B649B649B649B649B649B64DB24DB24D926D936C93649B64DB26D936C9B64DB26D936C9B24D936C9B64D936C9B24D93649B26C9B64D9364DB26C9B26C9B26D9364D9364D9364D9364D9364D9326C9B26C9B26CD9364D9326C9B264D9366C9B264D9326C99364C9B264D9B264D9326CD9326CD9B264D9B264C9B366C99326CD9B366C993264C9B366CD9B366CD9B366CD9B366CC993264C99B366CD993264CD9B3264CD9B3264CD993266CC99B3664CD9933664";

cyclonev_ram_block ram_block1a10(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "rom";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "clock0";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 8191;
defparam ram_block1a10.port_a_logical_ram_depth = 65536;
defparam ram_block1a10.port_a_logical_ram_width = 24;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init3 = "4CD9933664CD9B3266CC9933664C99B3664C99B3664C993366CD9B3264C993266CD9B366CD9B366CD9B366CD9B264C99326CD9B366C99326CD9B264C9B364C9B366C99366C99364C9B364C9B264D9326C99364C9B26CD9364C9B26C99364D9366C9B26C9B26C99364D9364D9364D9364D9364D936C9B26C9B26C9B64D9364DB26C9B24D93649B26D9364DB26D93649B26D936C9B64DB26D936C9B64DB24D926D936C93649B649B64DB24DB24DB24DB24DB24DB24DB24DB249B649B64936C936D926DB24DB649B6C926DB24DB64936D924DB64936DB249B6C924DB64926DB24936DB24936DB24926DB64924DB6C9249B6DB64924DB6DB24924DB6DB249249B6DB";
defparam ram_block1a10.mem_init2 = "6C924924DB6DB6D924924926DB6DB6DB64924924924936DB6DB6DB6DB6DB6C92492492492492492492492492492492492492492492DB6DB6DB6DB6DB6DA492492492492DB6DB6DB6924924925B6DB6DA4924925B6DB6D24924B6DB6D24924B6DB692492DB6DA4924B6DB4924B6DB4924B6DB4924B6DA4925B6D2496DB4925B6D2496DB4925B6D24B6DA496DB492DB6925B6925B6D24B6D24B6D24B6D24B6D24B6D25B6925B692DB492DA496DA4B6D25B692DB496DA4B6925B496DA4B6925B496D24B692DA4B6925B496D25B496D25B496D25B496D25B496D25B49692DA4B692DA5B496D25A4B692DA5B49692DA4B496D2DA4B496D2DA4B49692DA5B4B696D25A";
defparam ram_block1a10.mem_init1 = "4B49692D25A4B49692D25A4B49692D25A5B4B696D2D25A4B4B696D2D25A5B4B49696D2D25A5B4B49696D2D2DA5A4B4B4969692D2D25A5A4B4B4969696D2D2D25A5A5B4B4B4B6969696D2D2D2D25A5A5A5A4B4B4B4B4969696969692D2D2D2D2D2D2D25A5A5A5A5A5A5A5A5A5A5B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B5A5A5A5A5A5A5A5A5A5A5A5AD2D2D2D2D2D2D2969696969696B4B4B4B4B5A5A5A5A5AD2D2D2D296969694B4B4B4A5A5A5AD2D2D2969696B4B4B5A5A5A52D2D2969694B4B4A5A5AD2D2D69694B4B5A5A5AD2D29696B4B4A5A52D2D69694B4B5A5AD2D29694B4B5A5AD2D69694B4A5A52D29694B4A5A52D29694B4A5A52D29694";
defparam ram_block1a10.mem_init0 = "B4A5A52D696B4B5A52D29694B5A5AD2D694B4A5AD2D694B4A5AD2D694B5A5AD29694B5A52D296B4A5AD2D694B5A52D296B4A5AD29694B5A52D694B5A52D696B4A5AD296B4A5AD296B4A5AD296B4A5AD296B4A5AD296B4A52D694B5A52D694B5A5296B4A5AD296B4A52D694B5A5296B4A5AD294B5A52D6B4A5AD294B5A52D6B4A5AD294B5A5296B4A5AD694B5AD296B5A52D6B4A5AD694B5AD296B5A52D6B4A52D694A5AD294B5AD296B5A5296B4A52D6B4A5AD694A5AD294B5AD294B5A5296B5A5296B5A52D6B4A52D6B4A52D694A5AD694A5AD694A5AD694B5AD294B5AD294B5AD294B5AD294B5A5296B5A5296B5A5296B5A5296B5A5296B5A5296B5A5296B4";

cyclonev_ram_block ram_block1a34(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a34_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a34.clk0_core_clock_enable = "ena0";
defparam ram_block1a34.clk0_input_clock_enable = "ena0";
defparam ram_block1a34.clk0_output_clock_enable = "ena0";
defparam ram_block1a34.data_interleave_offset_in_bits = 1;
defparam ram_block1a34.data_interleave_width_in_bits = 1;
defparam ram_block1a34.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a34.init_file_layout = "port_a";
defparam ram_block1a34.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a34.operation_mode = "rom";
defparam ram_block1a34.port_a_address_clear = "none";
defparam ram_block1a34.port_a_address_width = 13;
defparam ram_block1a34.port_a_data_out_clear = "none";
defparam ram_block1a34.port_a_data_out_clock = "clock0";
defparam ram_block1a34.port_a_data_width = 1;
defparam ram_block1a34.port_a_first_address = 8192;
defparam ram_block1a34.port_a_first_bit_number = 10;
defparam ram_block1a34.port_a_last_address = 16383;
defparam ram_block1a34.port_a_logical_ram_depth = 65536;
defparam ram_block1a34.port_a_logical_ram_width = 24;
defparam ram_block1a34.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.ram_block_type = "auto";
defparam ram_block1a34.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFC00000000007FFFFFFFFF000000001FFFFFFFE0000000FFFFFFF0000001FFFFFF000000FFFFFE000007FFFFE00001FFFFF00001FFFFC0000FFFFC0000FFFF80003FFFE0001FFFE0003FFF8000FFFE0003FFF0003FFF0003FFE0007FFC001FFE000FFF8007FF8007FF8007FF800FFF001FFE003FF800FFE007FF001FF800FFC00FFC00FFC00FFC00FFC01FF801FF007FE00FF803FE007FC03FE00FF803FC01FF00FF807FC03FC03FE01FE01FE01FE01FE01FE01FC03FC03F807F00FE01FC03F807F01FE03F80FE03FC07F01FC07F01FC0FE03F80FC07F01F80FE07F03F8";
defparam ram_block1a34.mem_init2 = "1FC0FE07F03F01F80FC0FC07E07E07F03F03F03F03F03F03F03F03F03F03F07E07E07C0FC0F81F83F03E07C0FC1F83F07E0FC1F83F07C0F81F07E0F83F07C0F83E07C1F07C0F83E0F83E07C1F07C1F07C1F07C1F0783E0F83E0F87C1F07C3E0F87C1F0F83E1F0783E1F0783E1F0F83C1E0F07C3E1F0F87C3E1F0F0783C1E1F0F8783C3E1F0F0F8783C3E1E1F0F0F8787C3C3C1E1E1E0F0F0F0F878787878783C3C3C3C3C3C3C3C3C3C3C3C3C3C3C787878787870F0F0F1E1E1E1C3C3C787870F0F1E1E3C3C7878F0E1E1C3C7870F1E1C3C7870E1E3C3870F1E3C3870E1C3C78F1E3C78F1E3C78F1E3C78F1E3C78E1C3871E3C78E1C38F1C3871E3870E3C70E3C";
defparam ram_block1a34.mem_init1 = "70E3871E3871E38F1C78E1C70E3871C78E3C71E38E1C71E38E3C71C78E38F1C71C38E38E1C71C71E38E38E3871C71C71C71C38E38E38E38E38E38E38E38E38E38E38E38E39C71C71C71C718E38E38E31C71C738E38E31C71C638E39C71CE38E71C738E39C718E39C718E39C718E31C638E71CE39C738E718E31C639C738C718E718E31CE31CE31CE31CE31CE31CE31CE318E718C738C639C631CE718C739C6318E739C6318E739C6318C739CE739C6318C6318C6318E739CE739CE7318C6318C6318C6739CE7398C6318CE7398C6319CE7318CE7398C67398C67398C67398CE7319CE6339CC67318CE63398CE6319CC67319CC663398CE63398CC673198CE633";
defparam ram_block1a34.mem_init0 = "19CCE63319CCE673198CC663399CCE673399CCE6633198CC66733998CC66733998CCE66333998CCE66333199CCCE663331998CCC6663331999CCCE66633339998CCCC6666333319998CCCCE66663333399999CCCCCC6666673333339999999CCCCCCCE66666666333333333319999999999998CCCCCCCCCCCCCCCCCCCCCCCCCC666666666666666CCCCCCCCCCCCCCCCCCCCCCCCCC9999999999999B3333333333666666666CCCCCCCD999999B333333666666CCCCCD999993333366666CCCCD9999B33326666CCCC999933326664CCC99993336666CCC999B332666CCC999333666CCC999332664CC999332664CC99933666CC99933666CC99B33664CD993366";

cyclonev_ram_block ram_block1a107(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a107_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a107.clk0_core_clock_enable = "ena0";
defparam ram_block1a107.clk0_input_clock_enable = "ena0";
defparam ram_block1a107.clk0_output_clock_enable = "ena0";
defparam ram_block1a107.data_interleave_offset_in_bits = 1;
defparam ram_block1a107.data_interleave_width_in_bits = 1;
defparam ram_block1a107.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a107.init_file_layout = "port_a";
defparam ram_block1a107.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a107.operation_mode = "rom";
defparam ram_block1a107.port_a_address_clear = "none";
defparam ram_block1a107.port_a_address_width = 13;
defparam ram_block1a107.port_a_data_out_clear = "none";
defparam ram_block1a107.port_a_data_out_clock = "clock0";
defparam ram_block1a107.port_a_data_width = 1;
defparam ram_block1a107.port_a_first_address = 32768;
defparam ram_block1a107.port_a_first_bit_number = 11;
defparam ram_block1a107.port_a_last_address = 40959;
defparam ram_block1a107.port_a_logical_ram_depth = 65536;
defparam ram_block1a107.port_a_logical_ram_width = 24;
defparam ram_block1a107.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a107.ram_block_type = "auto";
defparam ram_block1a107.mem_init3 = "8F1E1C3878F1E3C3870F1E3C7870E1C3878F1E3C7870E1C3870E1C3C78F1E3C78F1E3C78F1E3C78F1E3C78F1E3C78F1E3C70E1C3870E1C38F1E3C78F1C3870E3C78F1E3870E1C78F1C3870E3C78E1C38F1E3870E3C70E1C78F1C38F1E3871E3870E3C70E3C70E1C78E1C78E1C78E1C78E1C78E1C70E3C70E3C70E3871E3871C38F1C38E1C78E3C71E3871C38E1C78E3C71E38F1C78E3C71E38F1C78E3C71E38E1C70E3871C78E3871C38E3C71C38E3C71C38E3C71C38E3C71C78E3871C70E38E1C71C38E3871C70E38E3C71C78E38E1C71C78E38E3C71C70E38E3871C71C38E38E3C71C71C38E38E3871C71C70E38E38E3871C71C71C38E38E38E3C71C71C71C";
defparam ram_block1a107.mem_init2 = "70E38E38E38E38E1C71C71C71C71C71C78E38E38E38E38E38E38E38E38E38F1C71C71C71C71C71C71C71C71C71C71C71C71C71C71CE38E38E38E38E38E38E38E38E38E31C71C71C71C71C71C638E38E38E38E39C71C71C71C738E38E38E38C71C71C71CE38E38E38C71C71C738E38E38C71C71C738E38E39C71C718E38E39C71C718E38E39C71C738E38E71C71CE38E39C71C638E38C71C738E38C71C738E38C71C638E39C71CE38E31C718E38C71C638E31C718E38C71C638E71C738E39C718E38C71CE38C71C638E71C638E71C638E71C638E71C638E71C638E71CE38C71CE39C718E39C738E31C638E71CE38C718E31C738E71CE38C718E31C638C718E39C";
defparam ram_block1a107.mem_init1 = "738E71CE39C738E71CE39C738E71CE39C638C718E31C638C738E71CE39C638C718E71CE39C638C718E71CE31C638C738E718E31CE39C638C738E718E71CE31C639C638C738C718E718E31CE31C639C639C738C738C718E718E718E31CE31CE31CE31C639C639C639C639C639C638C738C738C738C738C738C738C738C738C738C639C639C639C639C639C639CE31CE31CE31CE318E718E718E738C738C739C639C639CE31CE31CE718E718C738C739C639CE31CE318E718C738C639C639CE31CE718E738C739C631CE318E718C739C639CE31CE718C738C639CE318E718C739C631CE318E738C639CE318E718C739C631CE718C739C631CE718C739C631CE718";
defparam ram_block1a107.mem_init0 = "C739CE318E738C639CE318E739C631CE718C739CE318E738C631CE718C639CE318E739C631CE738C631CE718C639CE318C739CE318E739C6318E739C6318E738C631CE738C631CE738C631CE738C631CE738C631CE738C6318E739C6318E739C6318C739CE318C739CE718C639CE738C631CE739C6318C739CE318C639CE738C631CE739C6318C739CE718C631CE739C6318C739CE718C631CE739C6318C739CE718C631CE739CE318C639CE738C6318C739CE718C631CE739CE318C639CE739C6318C639CE738C6318C739CE718C6318E739CE718C6318E739CE318C631CE739CE318C631CE739C6318C639CE739C6318C639CE739C6318C639CE739C6318C6";

cyclonev_ram_block ram_block1a131(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a131_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a131.clk0_core_clock_enable = "ena0";
defparam ram_block1a131.clk0_input_clock_enable = "ena0";
defparam ram_block1a131.clk0_output_clock_enable = "ena0";
defparam ram_block1a131.data_interleave_offset_in_bits = 1;
defparam ram_block1a131.data_interleave_width_in_bits = 1;
defparam ram_block1a131.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a131.init_file_layout = "port_a";
defparam ram_block1a131.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a131.operation_mode = "rom";
defparam ram_block1a131.port_a_address_clear = "none";
defparam ram_block1a131.port_a_address_width = 13;
defparam ram_block1a131.port_a_data_out_clear = "none";
defparam ram_block1a131.port_a_data_out_clock = "clock0";
defparam ram_block1a131.port_a_data_width = 1;
defparam ram_block1a131.port_a_first_address = 40960;
defparam ram_block1a131.port_a_first_bit_number = 11;
defparam ram_block1a131.port_a_last_address = 49151;
defparam ram_block1a131.port_a_logical_ram_depth = 65536;
defparam ram_block1a131.port_a_logical_ram_width = 24;
defparam ram_block1a131.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a131.ram_block_type = "auto";
defparam ram_block1a131.mem_init3 = "0000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF8000000000000000001FFFFFFFFFFFFFFF00000000000001FFFFFFFFFFFF000000000007FFFFFFFFFE0000000001FFFFFFFFF000000000FFFFFFFFC00000001FFFFFFFC0000000FFFFFFFC0000003FFFFFFC0000007FFFFFE000000FFFFFF8000007FFFFF800000FFFFFE000003FFFFF000007FFFFE00000FFFFF00000FFFFF00000FFFFE00001FFFF80000FFFFC00007FFFC0000FFFFC0001FFFF00007FFFC0003FFFE0001FFFE0001FFFE0001FFFC0003FFF8000FFFE0003FFF8001FFFC000FFFC0007FFE0007FFE000FFFC000FFF8001FFF0007FFC00";
defparam ram_block1a131.mem_init2 = "1FFF0007FFC001FFF000FFF8007FF8003FFC003FFC003FFC003FFC003FFC007FF8007FF000FFE003FFC007FF001FFC007FF001FFC007FF003FF800FFC007FF003FF801FF800FFC00FFC007FE007FE007FE007FE007FC00FFC00FF801FF803FF007FE00FFC01FF803FE007FC01FF003FE00FF803FE00FF803FE00FF803FE01FF007FC03FE00FF007FC03FE01FF00FF807FC03FE01FE00FF00FF007F807F807FC03FC03FC03FC03FC03FC03FC03FC07F807F807F80FF00FE01FE01FC03F807F80FF01FE03FC07F80FF01FE03F807F01FE03F807F01FC03F80FE03FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07E03F80FE03F01FC07E03F80FC07F03F";
defparam ram_block1a131.mem_init1 = "80FC07E03F81FC0FE07F01F80FC07E07F03F81FC0FE07E03F03F81F80FC0FE07E03F03F01F81F81FC0FC0FC07E07E07E07E03F03F03F03F03F03F03F03F03F03F03F03F03E07E07E07E07E0FC0FC0FC1F81F83F03F03E07E07C0FC1F81F03F07E07C0FC1F81F03E07E0FC1F81F03E07C0F81F03E07C0F81F03E07C1F83F07E0F81F03E0FC1F03E0FC1F03E0FC1F03E0FC1F07E0F83F07C1F83E0F81F07C1F83E0F83E07C1F07C1F83E0F83E0F83E07C1F07C1F07C1F07C1F07C1F07C1F07C1F07C1F0783E0F83E0F83E0F07C1F07C1E0F83E0F07C1F0783E0F87C1F0783E0F07C1E0F83C1F0783E0F07C3E0F07C1E0F87C1E0F87C3E0F07C3E0F0783E1F0F83C";
defparam ram_block1a131.mem_init0 = "1E0F07C3E1F0F87C1E0F0783C1E0F0783C1E0F0783C1E0F0787C3E1F0F8783C1E0F0F87C3C1E0F0F87C3C1E1F0F0783C3E1E0F0F8783C3E1E1F0F0787C3C3E1E0F0F078783C3C1E1E0F0F0F8787C3C3C1E1E1F0F0F07878783C3C3C1E1E1E1F0F0F0F0787878783C3C3C3C3C1E1E1E1E1E1E1F0F0F0F0F0F0F0F0F0F0F0F0F0F878787878787878F0F0F0F0F0F0F0F0F0F0F0F0F0E1E1E1E1E1E1E3C3C3C3C3C3878787878F0F0F0F1E1E1E1C3C3C3C787878F0F0F1E1E1E3C3C387878F0F0E1E1E3C3C387870F0F1E1E3C3C7878F0F1E1E3C387870F0E1E3C3C7870F0E1E3C3878F0F1E1C3C7870F1E1C3C7870F1E1C3878F0E1E3C7870F1E3C3878F1E1C387";

cyclonev_ram_block ram_block1a155(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a155_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a155.clk0_core_clock_enable = "ena0";
defparam ram_block1a155.clk0_input_clock_enable = "ena0";
defparam ram_block1a155.clk0_output_clock_enable = "ena0";
defparam ram_block1a155.data_interleave_offset_in_bits = 1;
defparam ram_block1a155.data_interleave_width_in_bits = 1;
defparam ram_block1a155.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a155.init_file_layout = "port_a";
defparam ram_block1a155.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a155.operation_mode = "rom";
defparam ram_block1a155.port_a_address_clear = "none";
defparam ram_block1a155.port_a_address_width = 13;
defparam ram_block1a155.port_a_data_out_clear = "none";
defparam ram_block1a155.port_a_data_out_clock = "clock0";
defparam ram_block1a155.port_a_data_width = 1;
defparam ram_block1a155.port_a_first_address = 49152;
defparam ram_block1a155.port_a_first_bit_number = 11;
defparam ram_block1a155.port_a_last_address = 57343;
defparam ram_block1a155.port_a_logical_ram_depth = 65536;
defparam ram_block1a155.port_a_logical_ram_width = 24;
defparam ram_block1a155.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a155.ram_block_type = "auto";
defparam ram_block1a155.mem_init3 = "C3870F1E3C3878F1E1C3C78F0E1E3C3870F1E1C3C7870F1E1C3C7870F1E1E3C3878F0E1E1C3C7878F0E1E1C3C3878F0F1E1E3C3C7878F0F1E1E1C3C387878F0F0E1E1E3C3C387878F0F0F1E1E1E3C3C3C78787870F0F0F1E1E1E1E3C3C3C3C387878787878F0F0F0F0F0F0E1E1E1E1E1E1E1E1E1E1E1E1E1E3C3C3C3C3C3C3C3E1E1E1E1E1E1E1E1E1E1E1E1E1F0F0F0F0F0F0F078787878783C3C3C3C1E1E1E1F0F0F0F07878783C3C3C1E1E1F0F0F078787C3C3E1E1E0F0F078783C3C1E1E0F0F8787C3C1E1F0F0F8783C3E1E0F0F8783C1E1F0F0787C3E1E0F0787C3E1E0F0783C3E1F0F87C3C1E0F0783C1E0F0783C1E0F0783C1E0F07C3E1F0F87C1E0F0";
defparam ram_block1a155.mem_init2 = "783E1F0F83C1E0F87C1E0F87C3E0F07C3E0F07C1E0F87C1E0F83C1F0783E0F07C1E0F83C1F07C3E0F83C1F07C1E0F83E0F07C1F07C1E0F83E0F83E0F83C1F07C1F07C1F07C1F07C1F07C1F07C1F07C1F07C0F83E0F83E0F83F07C1F07C0F83E0F83F07C1F03E0F83F07C1F83E0FC1F07E0F81F07E0F81F07E0F81F07E0F81F03E0FC1F83F07C0F81F03E07C0F81F03E07C0F81F03F07E0FC0F81F03F07E07C0FC1F81F03F07E07C0FC0F81F81F83F03F07E07E07E0FC0FC0FC0FC0F81F81F81F81F81F81F81F81F81F81F81F81F80FC0FC0FC0FC07E07E07F03F03F01F81F80FC0FE07E03F03F81F80FC0FE07F03F81FC0FC07E03F01FC0FE07F03F80FC07E03";
defparam ram_block1a155.mem_init1 = "F81FC07E03F80FC07F01F80FE03F80FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F80FE03F807F01FC03F80FF01FC03F80FF01FE03FC07F80FF01FE03FC03F807F00FF00FE01FE03FC03FC03FC07F807F807F807F807F807F807F807FC03FC03FC01FE01FE00FF00FF807FC03FE01FF00FF807FC01FE00FF807FC01FF00FF803FE00FF803FE00FF803FE00FF801FF007FC00FF803FF007FE00FFC01FF803FF003FE007FE007FC00FFC00FFC00FFC00FFC007FE007FE003FF003FF801FFC007FE003FF801FFC007FF001FFC007FF001FFC007FF800FFE001FFC003FFC007FF8007FF8007FF8007FF8007FF8003FFC003FFE001FFF0007FFC001FFF0";
defparam ram_block1a155.mem_init0 = "007FFC001FFF0003FFE0007FFE000FFFC000FFFC0007FFE0007FFF0003FFF8000FFFE0003FFF80007FFF0000FFFF0000FFFF0000FFFF80007FFFC0001FFFF00007FFFE00007FFFC00007FFFE00003FFFF00000FFFFE00001FFFFE00001FFFFE00000FFFFFC00001FFFFF800000FFFFFE000003FFFFFC000003FFFFFE000000FFFFFFC0000007FFFFFF80000007FFFFFFE00000007FFFFFFF000000007FFFFFFFE000000001FFFFFFFFF0000000000FFFFFFFFFFC00000000001FFFFFFFFFFFF00000000000001FFFFFFFFFFFFFFF0000000000000000003FFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a179(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a179_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a179.clk0_core_clock_enable = "ena0";
defparam ram_block1a179.clk0_input_clock_enable = "ena0";
defparam ram_block1a179.clk0_output_clock_enable = "ena0";
defparam ram_block1a179.data_interleave_offset_in_bits = 1;
defparam ram_block1a179.data_interleave_width_in_bits = 1;
defparam ram_block1a179.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a179.init_file_layout = "port_a";
defparam ram_block1a179.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a179.operation_mode = "rom";
defparam ram_block1a179.port_a_address_clear = "none";
defparam ram_block1a179.port_a_address_width = 13;
defparam ram_block1a179.port_a_data_out_clear = "none";
defparam ram_block1a179.port_a_data_out_clock = "clock0";
defparam ram_block1a179.port_a_data_width = 1;
defparam ram_block1a179.port_a_first_address = 57344;
defparam ram_block1a179.port_a_first_bit_number = 11;
defparam ram_block1a179.port_a_last_address = 65535;
defparam ram_block1a179.port_a_logical_ram_depth = 65536;
defparam ram_block1a179.port_a_logical_ram_width = 24;
defparam ram_block1a179.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a179.ram_block_type = "auto";
defparam ram_block1a179.mem_init3 = "C6318C739CE738C6318C739CE738C6318C739CE738C6318C739CE718C6318E739CE718C6318E739CE318C631CE739CE318C631CE739C6318C639CE738C6318C739CE738C6318E739CE718C631CE739C6318C639CE738C6318E739CE718C631CE739C6318C739CE718C631CE739C6318C739CE718C631CE739C6318C739CE718C639CE738C6318E739C6318C739CE718C639CE738C631CE739C6318E739C6318C739CE318C739CE318C639CE718C639CE718C639CE718C639CE718C639CE718C639CE318C739CE318C739CE318E739C6318E738C631CE718C639CE718C739CE318E738C631CE718C639CE318E739C631CE718C739CE318E738C639CE318E739C6";
defparam ram_block1a179.mem_init2 = "31CE718C739C631CE718C739C631CE718C739C631CE318E738C639CE318E718C739C631CE318E738C639C631CE718E738C739C631CE318E718C739C639CE31CE718E738C738C639C631CE318E718E738C739C639C631CE31CE718E718E738C738C739C639C639CE31CE31CE318E718E718E718E738C738C738C738C738C738C639C639C639C639C639C639C639C639C639C638C738C738C738C738C738C718E718E718E718E31CE31CE31C639C639C738C738C718E718E31CE31C639C638C738C718E71CE31CE39C638C738E718E31CE39C638C718E71CE31C638C738E71CE31C638C738E71CE39C638C718E31C638C738E71CE39C738E71CE39C738E71CE39C";
defparam ram_block1a179.mem_init1 = "738E31C638C718E31C638E71CE39C718E31C638E71CE38C718E39C738E31C738E71C638E71CE38C71CE38C71CE38C71CE38C71CE38C71CE38C71C638E71C638E31C738E39C71CE38C71C638E31C718E38C71C638E31C718E38E71C738E38C71C638E39C71C638E39C71C638E38C71C738E38E71C71CE38E39C71C738E38E31C71C738E38E31C71C738E38E39C71C71C638E38E39C71C71C638E38E38E71C71C71C638E38E38E39C71C71C71C738E38E38E38E38C71C71C71C71C71C718E38E38E38E38E38E38E38E38E38E71C71C71C71C71C71C71C71C71C71C71C71C71C71C71E38E38E38E38E38E38E38E38E38E3C71C71C71C71C71C70E38E38E38E38E1C";
defparam ram_block1a179.mem_init0 = "71C71C71C78E38E38E3871C71C71C38E38E38E1C71C71C38E38E3871C71C78E38E3871C71C38E38E1C71C78E38E3C71C70E38E3C71C78E38E1C71C38E3871C70E38E1C71C38E3C71C78E3871C78E3871C78E3871C78E3871C38E3C71C38E1C70E38F1C78E3C71E38F1C78E3C71E38F1C78E3C70E3871C38F1C78E3C70E3871E3871C38F1C38E1C78E1C78E1C70E3C70E3C70E3C70E3C70E3C70E1C78E1C78E1C38F1C38F1E3871E3C70E1C78E1C38F1E3870E3C78E1C3871E3C70E1C38F1E3C78E1C3871E3C78F1E3870E1C3870E1C78F1E3C78F1E3C78F1E3C78F1E3C78F1E3C78F1E3C7870E1C3870E1C3C78F1E3C3870E1C3C78F1E1C3878F1E3C3870F1E3";

cyclonev_ram_block ram_block1a59(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a59_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a59.clk0_core_clock_enable = "ena0";
defparam ram_block1a59.clk0_input_clock_enable = "ena0";
defparam ram_block1a59.clk0_output_clock_enable = "ena0";
defparam ram_block1a59.data_interleave_offset_in_bits = 1;
defparam ram_block1a59.data_interleave_width_in_bits = 1;
defparam ram_block1a59.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a59.init_file_layout = "port_a";
defparam ram_block1a59.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a59.operation_mode = "rom";
defparam ram_block1a59.port_a_address_clear = "none";
defparam ram_block1a59.port_a_address_width = 13;
defparam ram_block1a59.port_a_data_out_clear = "none";
defparam ram_block1a59.port_a_data_out_clock = "clock0";
defparam ram_block1a59.port_a_data_width = 1;
defparam ram_block1a59.port_a_first_address = 16384;
defparam ram_block1a59.port_a_first_bit_number = 11;
defparam ram_block1a59.port_a_last_address = 24575;
defparam ram_block1a59.port_a_logical_ram_depth = 65536;
defparam ram_block1a59.port_a_logical_ram_width = 24;
defparam ram_block1a59.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a59.ram_block_type = "auto";
defparam ram_block1a59.mem_init3 = "3C78F0E1C3C7870E1E3C3870F1E1C3C78F0E1E3C3878F0E1E3C3878F0E1E1C3C7870F1E1E3C387870F1E1E3C3C7870F0E1E1C3C387870F0E1E1E3C3C787870F0F1E1E1C3C3C787870F0F0E1E1E1C3C3C38787878F0F0F0E1E1E1E1C3C3C3C3C787878787870F0F0F0F0F0F1E1E1E1E1E1E1E1E1E1E1E1E1E1C3C3C3C3C3C3C3C1E1E1E1E1E1E1E1E1E1E1E1E1E0F0F0F0F0F0F0F8787878787C3C3C3C3E1E1E1E0F0F0F0F878787C3C3C3E1E1E0F0F0F878783C3C1E1E1F0F0F8787C3C3E1E1F0F078783C3E1E0F0F0787C3C1E1F0F0787C3E1E0F0F8783C1E1F0F8783C1E1F0F87C3C1E0F0783C3E1F0F87C3E1F0F87C3E1F0F87C3E1F0F83C1E0F0783E1F0F";
defparam ram_block1a59.mem_init2 = "87C1E0F07C3E1F0783E1F0783C1F0F83C1F0F83E1F0783E1F07C3E0F87C1F0F83E1F07C3E0F83C1F07C3E0F83E1F07C1F0F83E0F83E1F07C1F07C1F07C3E0F83E0F83E0F83E0F83E0F83E0F83E0F83E0F83F07C1F07C1F07C0F83E0F83F07C1F07C0F83E0FC1F07C0F83E07C1F03E0F81F07E0F81F07E0F81F07E0F81F07E0FC1F03E07C0F83F07E0FC1F83F07E0FC1F83F07E0FC0F81F03F07E0FC0F81F83F03E07E0FC0F81F83F03F07E07E07C0FC0F81F81F81F03F03F03F03F07E07E07E07E07E07E07E07E07E07E07E07E07F03F03F03F03F81F81F80FC0FC0FE07E07F03F01F81FC0FC07E07F03F01F80FC07E03F03F81FC0FE03F01F80FC07F03F81FC";
defparam ram_block1a59.mem_init1 = "07E03F81FC07F03F80FE07F01FC07F03F80FE03F80FE03F80FE03F80FE03F80FE03F80FE03F807F01FC07F80FE03FC07F00FE03FC07F00FE01FC03F807F00FE01FC03FC07F80FF00FF01FE01FC03FC03FC03F807F807F807F807F807F807F807F803FC03FC03FE01FE01FF00FF007F803FC01FE00FF007F803FE01FF007F803FE00FF007FC01FF007FC01FF007FC01FF007FE00FF803FF007FC00FF801FF003FE007FC00FFC01FF801FF803FF003FF003FF003FF003FF801FF801FFC00FFC007FE003FF801FFC00FFE003FF800FFE003FF800FFE003FF8007FF001FFE003FFC003FF8007FF8007FF8007FF8007FF8007FFC003FFC001FFE000FFF8003FFE000F";
defparam ram_block1a59.mem_init0 = "FF8003FFE000FFFC001FFF8001FFF0003FFF0003FFF8001FFF8000FFFC0007FFF0001FFFC0007FFF8000FFFF0000FFFF0000FFFF00007FFF80003FFFE0000FFFF80001FFFF80003FFFF80001FFFFC0000FFFFF00001FFFFE00001FFFFE00001FFFFF000003FFFFE000007FFFFF000001FFFFFC000003FFFFFC000001FFFFFF0000003FFFFFF80000007FFFFFF80000001FFFFFFF80000000FFFFFFFF800000001FFFFFFFFE000000000FFFFFFFFFF00000000003FFFFFFFFFFE000000000000FFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFFFFFC000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a83(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a83_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a83.clk0_core_clock_enable = "ena0";
defparam ram_block1a83.clk0_input_clock_enable = "ena0";
defparam ram_block1a83.clk0_output_clock_enable = "ena0";
defparam ram_block1a83.data_interleave_offset_in_bits = 1;
defparam ram_block1a83.data_interleave_width_in_bits = 1;
defparam ram_block1a83.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a83.init_file_layout = "port_a";
defparam ram_block1a83.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a83.operation_mode = "rom";
defparam ram_block1a83.port_a_address_clear = "none";
defparam ram_block1a83.port_a_address_width = 13;
defparam ram_block1a83.port_a_data_out_clear = "none";
defparam ram_block1a83.port_a_data_out_clock = "clock0";
defparam ram_block1a83.port_a_data_width = 1;
defparam ram_block1a83.port_a_first_address = 24576;
defparam ram_block1a83.port_a_first_bit_number = 11;
defparam ram_block1a83.port_a_last_address = 32767;
defparam ram_block1a83.port_a_logical_ram_depth = 65536;
defparam ram_block1a83.port_a_logical_ram_width = 24;
defparam ram_block1a83.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a83.ram_block_type = "auto";
defparam ram_block1a83.mem_init3 = "39CE738C6318C739CE738C6318C739CE738C6318C739CE738C6318E739CE718C6318E739CE718C631CE739CE318C631CE739CE318C639CE739C6318C739CE738C6318C739CE718C6318E739CE318C639CE739C6318C739CE718C6318E739CE318C639CE738C6318E739CE318C639CE738C6318E739CE318C639CE738C6318E739C6318C739CE718C639CE738C6318E739C6318C739CE318C639CE718C639CE738C631CE738C631CE739C6318E739C6318E739C6318E739C6318E739C6318E739C631CE738C631CE738C631CE718C639CE718C739CE318E739C6318E738C631CE718C739CE318E739C631CE718C639CE318E738C631CE718C739C631CE738C639";
defparam ram_block1a83.mem_init2 = "CE318E738C639CE318E738C639CE318E738C639CE31CE718C739C631CE718E738C639CE31CE718C739C639CE318E718C738C639CE31CE718E738C639C631CE318E718C738C739C639CE31CE718E718C738C639C639CE31CE318E718E718C738C738C639C639C631CE31CE31CE718E718E718E718C738C738C738C738C738C739C639C639C639C639C639C639C639C639C639C738C738C738C738C738C738E718E718E718E71CE31CE31CE39C639C638C738C738E718E71CE31CE39C639C738C738E718E31CE31C639C738C718E71CE31C639C738E718E31CE39C738C718E31CE39C738C718E31C639C738E71CE39C738C718E31C638C718E31C638C718E31C63";
defparam ram_block1a83.mem_init1 = "8C71CE39C738E71CE39C718E31C638E71CE39C718E31C738E71C638C71CE38C718E39C718E31C738E31C738E31C738E31C738E31C738E31C738E39C718E39C71CE38C71C638E31C738E39C71CE38E71C738E39C71CE38E71C718E38C71C738E39C71C638E39C71C638E39C71C738E38C71C718E38E31C71C638E38C71C71CE38E38C71C71CE38E38C71C71C638E38E39C71C71C638E38E39C71C71C718E38E38E39C71C71C71C638E38E38E38C71C71C71C71C738E38E38E38E38E38E71C71C71C71C71C71C71C71C71C718E38E38E38E38E38E38E38E38E38E38E38E38E38E38E1C71C71C71C71C71C71C71C71C71C38E38E38E38E38E38F1C71C71C71C71E3";
defparam ram_block1a83.mem_init0 = "8E38E38E3871C71C71C78E38E38E3C71C71C71E38E38E3C71C71C78E38E3871C71C78E38E3C71C71E38E3871C71C38E38F1C71C38E3871C71E38E3C71C78E38F1C71E38E3C71C38E3871C78E3871C78E3871C78E3871C78E3C71C38E3C71E38F1C70E3871C38E1C70E3871C38E1C70E3871C38F1C78E3C70E3871C38F1C78E1C78E3C70E3C71E3871E3871E38F1C38F1C38F1C38F1C38F1C38F1E3871E3871E3C70E3C70E1C78E1C38F1E3871E3C70E1C78F1C3871E3C78E1C38F1E3C70E1C3871E3C78E1C3870E1C78F1E3C78F1E3870E1C3870E1C3870E1C3870E1C3870E1C3870E1C3878F1E3C78F1E3C3870E1C3C78F1E3C3870E1E3C7870E1C3C78F0E1C";

cyclonev_ram_block ram_block1a11(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "rom";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "clock0";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 8191;
defparam ram_block1a11.port_a_logical_ram_depth = 65536;
defparam ram_block1a11.port_a_logical_ram_width = 24;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init3 = "70E1E3C7870E1C3C78F0E1C3878F1E3C7870E1C3878F1E3C78F1E3C3870E1C3870E1C3870E1C3870E1C3870E1C3870E1C38F1E3C78F1E3C70E1C3870E3C78F1C3870E1C78F1E3870E3C78F1C3871E3C70E1C78F1C38F1E3870E3C70E1C78E1C78F1C38F1C38F1E3871E3871E3871E3871E3871E38F1C38F1C38F1C78E1C78E3C70E3C71E3871C38E1C78E3C71E3871C38E1C70E3871C38E1C70E3871C38E1C71E38F1C78E3871C78E3C71C38E3C71C38E3C71C38E3C71C38E3871C78E38F1C71E38E3C71C78E38F1C71C38E3871C71E38E3871C71C38E38F1C71C78E38E3C71C71C38E38E3C71C71C78E38E38F1C71C71C78E38E38E3C71C71C71C38E38E38E3";
defparam ram_block1a11.mem_init2 = "8F1C71C71C71C71E38E38E38E38E38E3871C71C71C71C71C71C71C71C71C70E38E38E38E38E38E38E38E38E38E38E38E38E38E38E31C71C71C71C71C71C71C71C71C71CE38E38E38E38E38E39C71C71C71C71C638E38E38E38C71C71C71C738E38E38E31C71C71C738E38E38C71C71C738E38E38C71C71C638E38E71C71C638E38E71C71C638E38C71C718E38E31C71C638E39C71C738E38C71C738E38C71C738E39C71C638E31C71CE38E71C738E39C71CE38E71C738E39C718E38C71C638E71C738E31C738E39C718E39C718E39C718E39C718E39C718E39C718E31C738E31C638E71C638C71CE39C718E31C738E71CE38C718E31C738E71CE39C738E71C63";
defparam ram_block1a11.mem_init1 = "8C718E31C638C718E31C638C718E31C639C738E71CE39C738C718E31C639C738E718E31C639C738E718E31CE39C738C718E71CE31C639C738C718E718E31CE39C639C738C738E718E71CE31CE39C639C638C738C738E718E718E71CE31CE31CE31CE39C639C639C639C639C639C738C738C738C738C738C738C738C738C738C739C639C639C639C639C639C631CE31CE31CE31CE718E718E718C738C738C639C639C631CE31CE318E718E738C738C639C631CE31CE718E738C739C639C631CE318E718C738C639CE31CE718E738C639C631CE318E738C739C631CE718E738C639CE31CE718C739C631CE718E738C639CE318E738C639CE318E738C639CE318E7";
defparam ram_block1a11.mem_init0 = "38C639CE718C739C631CE718C639CE318E738C631CE718C739CE318E739C631CE718C639CE318C739CE318E739C631CE738C631CE718C639CE718C639CE718C739CE318C739CE318C739CE318C739CE318C739CE318C739CE718C639CE718C639CE738C631CE738C6318E739C6318C739CE318C639CE738C631CE739C6318C739CE318C639CE738C6318E739CE318C639CE738C6318E739CE318C639CE738C6318E739CE318C631CE739C6318C739CE738C6318E739CE318C631CE739C6318C639CE739C6318C739CE738C6318E739CE718C6318E739CE718C631CE739CE318C631CE739CE318C639CE739C6318C639CE739C6318C639CE739C6318C639CE738";

cyclonev_ram_block ram_block1a35(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a35_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a35.clk0_core_clock_enable = "ena0";
defparam ram_block1a35.clk0_input_clock_enable = "ena0";
defparam ram_block1a35.clk0_output_clock_enable = "ena0";
defparam ram_block1a35.data_interleave_offset_in_bits = 1;
defparam ram_block1a35.data_interleave_width_in_bits = 1;
defparam ram_block1a35.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a35.init_file_layout = "port_a";
defparam ram_block1a35.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a35.operation_mode = "rom";
defparam ram_block1a35.port_a_address_clear = "none";
defparam ram_block1a35.port_a_address_width = 13;
defparam ram_block1a35.port_a_data_out_clear = "none";
defparam ram_block1a35.port_a_data_out_clock = "clock0";
defparam ram_block1a35.port_a_data_width = 1;
defparam ram_block1a35.port_a_first_address = 8192;
defparam ram_block1a35.port_a_first_bit_number = 11;
defparam ram_block1a35.port_a_last_address = 16383;
defparam ram_block1a35.port_a_logical_ram_depth = 65536;
defparam ram_block1a35.port_a_logical_ram_width = 24;
defparam ram_block1a35.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.ram_block_type = "auto";
defparam ram_block1a35.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000007FFFFFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFE000000000000FFFFFFFFFFF80000000001FFFFFFFFFE000000000FFFFFFFFF000000003FFFFFFFE00000003FFFFFFF00000003FFFFFFC0000003FFFFFF8000001FFFFFF0000007FFFFF8000007FFFFF000001FFFFFC00000FFFFF800001FFFFF00000FFFFF00000FFFFF00001FFFFE00007FFFF00003FFFF80003FFFF00003FFFE0000FFFF80003FFFC0001FFFE0001FFFE0001FFFE0003FFFC0007FFF0001FFFC0007FFE0003FFF0003FFF8001FFF8001FFF0003FFF0007FFE000FFF8003FF";
defparam ram_block1a35.mem_init2 = "E000FFF8003FFE000FFF0007FF8007FFC003FFC003FFC003FFC003FFC003FF8007FF800FFF001FFC003FF800FFE003FF800FFE003FF800FFE007FF003FF800FFC007FE007FF003FF003FF801FF801FF801FF801FF803FF003FF007FE007FC00FF801FF003FE007FC01FF803FE00FFC01FF007FC01FF007FC01FF007FC01FE00FF803FC01FF00FF803FC01FE00FF007F803FC01FE01FF00FF00FF807F807F803FC03FC03FC03FC03FC03FC03FC03F807F807F807F00FF01FE01FE03FC07F807F00FE01FC03F807F00FE01FC07F80FE01FC07F80FE03FC07F01FC03F80FE03F80FE03F80FE03F80FE03F80FE03F80FE03F81FC07F01FC0FE03F81FC07F03F80FC0";
defparam ram_block1a35.mem_init1 = "7F03F81FC07E03F01F80FE07F03F81F80FC07E03F01F81FC0FC07E07F03F01F81FC0FC0FE07E07E03F03F03F81F81F81F81FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC1F81F81F81F81F03F03F03E07E07C0FC0FC1F81F83F03E07E0FC0F81F83F03E07E0FC1F81F03E07E0FC1F83F07E0FC1F83F07E0FC1F83E07C0F81F07E0FC1F03E0FC1F03E0FC1F03E0FC1F03E0F81F07C0F83E07C1F07E0F83E07C1F07C1F83E0F83E07C1F07C1F07C1F83E0F83E0F83E0F83E0F83E0F83E0F83E0F83E0F87C1F07C1F07C1F0F83E0F83E1F07C1F0F83E0F87C1F0783E0F87C1F0F83E1F07C3E0F87C1F0F83C1F0F83E1F0783E1F0783C1F0F83C1F0F87C1E0F07C3";
defparam ram_block1a35.mem_init0 = "E1F0F83C1E0F0783E1F0F87C3E1F0F87C3E1F0F87C3E1F0F8783C1E0F0787C3E1F0F0783C3E1F0F0783C3E1E0F0F87C3C1E1F0F0787C3C1E1E0F0F8783C3C1E1F0F0F8787C3C3E1E1F0F0F078783C3C3E1E1E0F0F0F878787C3C3C3E1E1E1E0F0F0F0F87878787C3C3C3C3C3E1E1E1E1E1E1E0F0F0F0F0F0F0F0F0F0F0F0F0F07878787878787870F0F0F0F0F0F0F0F0F0F0F0F0F1E1E1E1E1E1E1C3C3C3C3C3C7878787870F0F0F0E1E1E1E3C3C3C38787870F0F0E1E1E1C3C3C787870F0F1E1E1C3C3C7878F0F0E1E1C3C387870F0E1E1C3C7878F0F1E1C3C3878F0F1E1C3C7870F0E1E3C3878F0E1E3C3878F0E1E3C7870F1E1C3878F0E1C3C7870E1E3C78";

cyclonev_ram_block ram_block1a108(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a108_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a108.clk0_core_clock_enable = "ena0";
defparam ram_block1a108.clk0_input_clock_enable = "ena0";
defparam ram_block1a108.clk0_output_clock_enable = "ena0";
defparam ram_block1a108.data_interleave_offset_in_bits = 1;
defparam ram_block1a108.data_interleave_width_in_bits = 1;
defparam ram_block1a108.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a108.init_file_layout = "port_a";
defparam ram_block1a108.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a108.operation_mode = "rom";
defparam ram_block1a108.port_a_address_clear = "none";
defparam ram_block1a108.port_a_address_width = 13;
defparam ram_block1a108.port_a_data_out_clear = "none";
defparam ram_block1a108.port_a_data_out_clock = "clock0";
defparam ram_block1a108.port_a_data_width = 1;
defparam ram_block1a108.port_a_first_address = 32768;
defparam ram_block1a108.port_a_first_bit_number = 12;
defparam ram_block1a108.port_a_last_address = 40959;
defparam ram_block1a108.port_a_logical_ram_depth = 65536;
defparam ram_block1a108.port_a_logical_ram_width = 24;
defparam ram_block1a108.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a108.ram_block_type = "auto";
defparam ram_block1a108.mem_init3 = "80FE03F807F01FC07F00FE03F80FE03F807F01FC07F01FC07F01FC03F80FE03F80FE03F80FE03F80FE03F80FE03F80FE03F01FC07F01FC07F01FC07F03F80FE03F80FE07F01FC07F03F80FE03F81FC07F01F80FE03F01FC07F03F80FE07F01F80FE03F01FC0FE03F81FC07E03F81FC07E03F81FC0FE03F01FC0FE07F01F80FC07F03F81FC07E03F01F80FC07E03F81FC0FE07F03F81FC0FE07F03F81FC0FE07E03F01F80FC07E07F03F81FC0FC07E03F03F81FC0FC07E03F03F81F80FC0FE07E03F03F81F80FC0FE07E03F03F81F81FC0FC07E07E03F03F01F81F80FC0FC07E07E03F03F03F81F81F80FC0FC0FE07E07E07F03F03F03F81F81F81FC0FC0FC0FC";
defparam ram_block1a108.mem_init2 = "0FE07E07E07E07E03F03F03F03F03F03F81F81F81F81F81F81F81F81F81F80FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC1F81F81F81F81F81F81F81F81F81F03F03F03F03F03F03E07E07E07E07E07C0FC0FC0FC0F81F81F81F83F03F03F03E07E07E07C0FC0FC0F81F81F83F03F03F07E07E07C0FC0F81F81F83F03F07E07E07C0FC0F81F81F03F03E07E07C0FC1F81F83F03F07E07C0FC0F81F83F03E07E07C0FC1F81F03F07E07C0FC1F81F03F07E07C0FC1F81F03F07E07C0F81F83F03E07C0FC1F81F03E07E0FC1F81F03E07E0FC1F81F03E07E0FC1F83F03E07C0F81F83F07E0FC1F81F03E07C0F81F03F07E0FC1F83F07E0FC1F83F07E07C";
defparam ram_block1a108.mem_init1 = "0F81F03E07C0F81F03E07C0F81F03E07C1F83F07E0FC1F83F07E0FC1F83E07C0F81F03E07C1F83F07E0FC1F03E07C0F81F07E0FC1F83E07C0F81F07E0FC1F03E07C1F83F07C0F81F07E0FC1F03E07C1F83F07C0F83F07E0F81F07E0FC1F03E0FC1F03E07C1F83E07C1F83E07C1F83F07C0F83F07C0F83F07C0F83F07C0F83F07C1F83E07C1F83E07C1F83E07C1F03E0FC1F03E0F81F07E0F81F07C0F83F07C1F83E07C1F03E0FC1F07E0F83F07C0F83E07C1F03E0F81F07C0F83E07C1F83E0FC1F07E0F83F07C1F03E0F81F07C0F83E07C1F03E0F83F07C1F83E0F81F07C0F83E0FC1F07E0F83E07C1F07E0F83F07C1F03E0F83F07C1F03E0F83F07C1F03E0F8";
defparam ram_block1a108.mem_init0 = "3F07C1F07E0F83E07C1F07E0F83E0FC1F07C0F83E0F81F07C1F03E0F83E07C1F07E0F83E0FC1F07C1F03E0F83E07C1F07C0F83E0F81F07C1F07E0F83E0F81F07C1F03E0F83E0FC1F07C1F03E0F83E0FC1F07C1F03E0F83E0F81F07C1F07E0F83E0F83F07C1F07C0F83E0F83E07C1F07C1F03E0F83E0F83F07C1F07C1F83E0F83E0FC1F07C1F07C0F83E0F83E0FC1F07C1F07C0F83E0F83E0FC1F07C1F07C0F83E0F83E0FC1F07C1F07C1F83E0F83E0F83F07C1F07C1F03E0F83E0F83E07C1F07C1F07C1F83E0F83E0F83F07C1F07C1F07E0F83E0F83E0F81F07C1F07C1F03E0F83E0F83E0FC1F07C1F07C1F83E0F83E0F83E07C1F07C1F07C1F83E0F83E0F83E";

cyclonev_ram_block ram_block1a132(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a132_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a132.clk0_core_clock_enable = "ena0";
defparam ram_block1a132.clk0_input_clock_enable = "ena0";
defparam ram_block1a132.clk0_output_clock_enable = "ena0";
defparam ram_block1a132.data_interleave_offset_in_bits = 1;
defparam ram_block1a132.data_interleave_width_in_bits = 1;
defparam ram_block1a132.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a132.init_file_layout = "port_a";
defparam ram_block1a132.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a132.operation_mode = "rom";
defparam ram_block1a132.port_a_address_clear = "none";
defparam ram_block1a132.port_a_address_width = 13;
defparam ram_block1a132.port_a_data_out_clear = "none";
defparam ram_block1a132.port_a_data_out_clock = "clock0";
defparam ram_block1a132.port_a_data_width = 1;
defparam ram_block1a132.port_a_first_address = 40960;
defparam ram_block1a132.port_a_first_bit_number = 12;
defparam ram_block1a132.port_a_last_address = 49151;
defparam ram_block1a132.port_a_logical_ram_depth = 65536;
defparam ram_block1a132.port_a_logical_ram_width = 24;
defparam ram_block1a132.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a132.ram_block_type = "auto";
defparam ram_block1a132.mem_init3 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFE0000000000000000000FFFFFFFFFFFFFFFFFC0000000000000003FFFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFE0000000000007FFFFFFFFFFF800000000001FFFFFFFFFFF00000000001FFFFFFFFFF0000000000FFFFFFFFFE0000000007FFFFFFFFC000000003FFFFFFFFC00000000FFFFFFFFC00000001FFFFFFFE00000001FFFFFFFC00000007FFFFFFE00000007FFFFFFC0000003FFFFFFE0000001FFFFFFC0000007FFFFFF0000003FF";
defparam ram_block1a132.mem_init2 = "FFFF0000003FFFFFF0000007FFFFF8000003FFFFFC000003FFFFFC000003FFFFF800000FFFFFE000003FFFFF000003FFFFF000003FFFFF000007FFFFC00000FFFFF800007FFFFC00003FFFFE00001FFFFE00001FFFFC00003FFFF800007FFFF00001FFFFC00007FFFE00003FFFF00001FFFF80001FFFF80001FFFF80001FFFF00003FFFE0000FFFFC0001FFFF00007FFFC0001FFFE0000FFFF00007FFF80003FFFC0003FFFC0003FFFC0003FFFC0007FFF80007FFF0001FFFE0003FFF80007FFF0001FFFC0007FFF0001FFF8000FFFE0007FFF0003FFF8001FFFC000FFFC000FFFC000FFFC000FFFC000FFFC000FFFC001FFF8001FFF0003FFE0007FFC000FFF";
defparam ram_block1a132.mem_init1 = "8003FFE0007FFC001FFF0007FFC001FFF0007FFC001FFE000FFF8007FFC001FFE000FFF0007FF8003FFC003FFE001FFE001FFF000FFF000FFF000FFF000FFF000FFF000FFE001FFE001FFE003FFC003FF8007FF000FFE001FFC003FF800FFF001FFC003FF800FFE001FFC007FF001FFC007FF001FFC007FF001FFC007FF001FF800FFE003FF001FFC00FFE003FF001FFC00FFE007FF003FF801FF800FFC007FE007FE003FF003FF801FF801FF801FFC00FFC00FFC00FFC00FFC00FFC00FFC00FFC00FF801FF801FF801FF003FF003FE007FE00FFC00FF801FF803FF007FE00FFC01FF803FF007FE00FFC01FF003FE007FC01FF803FE00FFC01FF007FE00FF803";
defparam ram_block1a132.mem_init0 = "FE00FFC01FF007FC01FF007FC01FF007FC01FF007FC01FF007FC01FF007F803FE00FF803FC01FF007FC03FE00FF007FC01FE00FF807FC01FE00FF007FC03FE01FF00FF807FC03FE01FF00FF807FC03FC01FE00FF00FF807F803FC03FE01FE00FF00FF007F807F803FC03FC03FE01FE01FE01FF00FF00FF00FF00FF00FF00FF007F807F807F807F80FF00FF00FF00FF00FF00FF00FE01FE01FE01FE03FC03FC03F807F807F80FF00FF01FE01FC03FC03F807F80FF00FE01FE03FC07F807F00FE01FE03FC07F80FF00FE01FC03F807F00FE01FC07F80FF01FE03FC07F00FE01FC07F80FF01FC03F80FF01FC03F80FF01FC07F80FE01FC07F00FE03F807F01FC07F";

cyclonev_ram_block ram_block1a156(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a156_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a156.clk0_core_clock_enable = "ena0";
defparam ram_block1a156.clk0_input_clock_enable = "ena0";
defparam ram_block1a156.clk0_output_clock_enable = "ena0";
defparam ram_block1a156.data_interleave_offset_in_bits = 1;
defparam ram_block1a156.data_interleave_width_in_bits = 1;
defparam ram_block1a156.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a156.init_file_layout = "port_a";
defparam ram_block1a156.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a156.operation_mode = "rom";
defparam ram_block1a156.port_a_address_clear = "none";
defparam ram_block1a156.port_a_address_width = 13;
defparam ram_block1a156.port_a_data_out_clear = "none";
defparam ram_block1a156.port_a_data_out_clock = "clock0";
defparam ram_block1a156.port_a_data_width = 1;
defparam ram_block1a156.port_a_first_address = 49152;
defparam ram_block1a156.port_a_first_bit_number = 12;
defparam ram_block1a156.port_a_last_address = 57343;
defparam ram_block1a156.port_a_logical_ram_depth = 65536;
defparam ram_block1a156.port_a_logical_ram_width = 24;
defparam ram_block1a156.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a156.ram_block_type = "auto";
defparam ram_block1a156.mem_init3 = "FC07F01FC03F80FE01FC07F00FE03FC07F01FE03F807F01FE03F807F01FE03FC07F00FE01FC07F80FF01FE03FC07F00FE01FC03F807F00FE01FE03FC07F80FF00FE01FC03FC07F80FF00FE01FE03FC03F807F807F00FF01FE01FE03FC03FC03F807F807F80FF00FF00FF00FE01FE01FE01FE01FE01FE01FE03FC03FC03FC03FC01FE01FE01FE01FE01FE01FE01FF00FF00FF00FF807F807F803FC03FC01FE01FE00FF00FF807F803FC03FE01FE00FF007F807FC03FE01FF00FF807FC03FE01FF00FF807FC01FE00FF007FC03FE00FF007FC01FE00FF807FC01FF007F803FE00FF803FC01FF007FC01FF007FC01FF007FC01FF007FC01FF007FC01FF007FE00FF";
defparam ram_block1a156.mem_init2 = "803FE00FFC01FF007FE00FF803FF007FC00FF801FF007FE00FFC01FF803FF007FE00FFC01FF803FF003FE007FE00FFC00FF801FF801FF003FF003FF003FE007FE007FE007FE007FE007FE007FE007FE007FF003FF003FF003FF801FF800FFC00FFC007FE003FF003FF801FFC00FFE007FF001FF800FFE007FF001FF800FFE003FF001FFC007FF001FFC007FF001FFC007FF001FFC007FF000FFE003FF8007FF001FFE003FF8007FF000FFE001FFC003FF8007FF800FFF000FFF000FFE001FFE001FFE001FFE001FFE001FFE001FFF000FFF000FFF8007FF8003FFC001FFE000FFF0007FFC003FFE000FFF0007FFC001FFF0007FFC001FFF0007FFC000FFF8003";
defparam ram_block1a156.mem_init1 = "FFE0007FFC000FFF8001FFF0003FFF0007FFE0007FFE0007FFE0007FFE0007FFE0007FFE0007FFF0003FFF8001FFFC000FFFE0003FFF0001FFFC0007FFF0001FFFC0003FFF8000FFFF0001FFFC0003FFFC0007FFF80007FFF80007FFF80007FFF80003FFFC0001FFFE0000FFFF00007FFFC0001FFFF00007FFFE0000FFFF80001FFFF00003FFFF00003FFFF00003FFFF00001FFFF80000FFFFC00007FFFF00001FFFFC00003FFFF800007FFFF00000FFFFF00000FFFFF800007FFFFC00003FFFFE000007FFFFC00001FFFFF800001FFFFF800001FFFFF800000FFFFFE000003FFFFF8000007FFFFF8000007FFFFF8000003FFFFFC000001FFFFFF8000001FFFF";
defparam ram_block1a156.mem_init0 = "FF8000001FFFFFFC0000007FFFFFF0000000FFFFFFF80000007FFFFFFC0000000FFFFFFFC00000007FFFFFFF00000000FFFFFFFF000000007FFFFFFFE000000007FFFFFFFF8000000007FFFFFFFFC000000000FFFFFFFFFE0000000001FFFFFFFFFF00000000001FFFFFFFFFFF000000000003FFFFFFFFFFFC000000000000FFFFFFFFFFFFF800000000000007FFFFFFFFFFFFFF80000000000000007FFFFFFFFFFFFFFFFE0000000000000000000FFFFFFFFFFFFFFFFFFFFFE00000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a180(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a180_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a180.clk0_core_clock_enable = "ena0";
defparam ram_block1a180.clk0_input_clock_enable = "ena0";
defparam ram_block1a180.clk0_output_clock_enable = "ena0";
defparam ram_block1a180.data_interleave_offset_in_bits = 1;
defparam ram_block1a180.data_interleave_width_in_bits = 1;
defparam ram_block1a180.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a180.init_file_layout = "port_a";
defparam ram_block1a180.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a180.operation_mode = "rom";
defparam ram_block1a180.port_a_address_clear = "none";
defparam ram_block1a180.port_a_address_width = 13;
defparam ram_block1a180.port_a_data_out_clear = "none";
defparam ram_block1a180.port_a_data_out_clock = "clock0";
defparam ram_block1a180.port_a_data_width = 1;
defparam ram_block1a180.port_a_first_address = 57344;
defparam ram_block1a180.port_a_first_bit_number = 12;
defparam ram_block1a180.port_a_last_address = 65535;
defparam ram_block1a180.port_a_logical_ram_depth = 65536;
defparam ram_block1a180.port_a_logical_ram_width = 24;
defparam ram_block1a180.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a180.ram_block_type = "auto";
defparam ram_block1a180.mem_init3 = "F83E0F83E0F83F07C1F07C1F07C0F83E0F83E0F83F07C1F07C1F07E0F83E0F83E0F81F07C1F07C1F03E0F83E0F83E0FC1F07C1F07C1F83E0F83E0F83F07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F83E0F83E0F83F07C1F07C1F07E0F83E0F83E07C1F07C1F07E0F83E0F83E07C1F07C1F07E0F83E0F83E07C1F07C1F07E0F83E0F83F07C1F07C1F83E0F83E0F81F07C1F07C0F83E0F83E07C1F07C1F83E0F83E0FC1F07C1F03E0F83E0F81F07C1F07E0F83E0F81F07C1F07E0F83E0F81F07C1F03E0F83E0FC1F07C1F03E0F83E07C1F07C0F83E0F81F07C1F07E0F83E0FC1F07C0F83E0F81F07C1F03E0F83E07C1F07E0F83E0FC1F07C0F83E0FC1F07C1F8";
defparam ram_block1a180.mem_init2 = "3E0F81F07C1F83E0F81F07C1F83E0F81F07C1F83E0FC1F07C0F83E0FC1F07E0F83E07C1F03E0F83F07C1F83E0F81F07C0F83E07C1F03E0F81F07C1F83E0FC1F07E0F83F07C0F83E07C1F03E0F81F07C0F83E07C1F83E0FC1F07E0F81F07C0F83F07C1F83E07C1F03E0FC1F03E0F81F07E0F81F07C0F83F07C0F83F07C0F83F07C1F83E07C1F83E07C1F83E07C1F83E07C1F83F07C0F83F07C0F83F07C0F81F07E0F81F07E0FC1F03E0FC1F83E07C1F83F07C0F81F07E0FC1F03E07C1F83F07C0F81F07E0FC1F03E07C0F83F07E0FC1F03E07C0F81F07E0FC1F83F07C0F81F03E07C0F83F07E0FC1F83F07E0FC1F83F07C0F81F03E07C0F81F03E07C0F81F03E0";
defparam ram_block1a180.mem_init1 = "7C0FC1F83F07E0FC1F83F07E0FC1F81F03E07C0F81F03F07E0FC1F83F03E07C0F81F83F07E0FC0F81F03F07E0FC0F81F03F07E0FC0F81F03F07E07C0F81F83F03E07C0FC1F81F03F07E07C0FC1F81F03F07E07C0FC1F81F03F07E07C0FC0F81F83F03E07E07C0FC1F81F83F03F07E07C0FC0F81F81F03F03E07E07C0FC0FC1F81F83F03F03E07E07C0FC0FC1F81F81F83F03F03E07E07E07C0FC0FC0F81F81F81F83F03F03F03E07E07E07E07C0FC0FC0FC0FC0F81F81F81F81F81F81F03F03F03F03F03F03F03F03F03F07E07E07E07E07E07E07E07E07E07E07E07E07E07E07E03F03F03F03F03F03F03F03F03F03F81F81F81F81F81F80FC0FC0FC0FC0FE0";
defparam ram_block1a180.mem_init0 = "7E07E07E07F03F03F03F81F81F81FC0FC0FC0FE07E07E03F03F03F81F81F80FC0FC07E07E03F03F01F81F80FC0FC07E07F03F03F81F80FC0FE07E03F03F81F80FC0FE07E03F03F81F80FC07E07F03F81F80FC07E07F03F81FC0FC07E03F01F80FC0FE07F03F81FC0FE07F03F81FC0FE07F03F80FC07E03F01F80FC07F03F81FC07E03F01FC0FE07F01F80FE07F03F80FC07F03F80FC07F03F80FE07F01F80FE03F01FC0FE03F81FC07F01F80FE03F01FC07F03F80FE03F81FC07F01FC0FE03F80FE03F81FC07F01FC07F01FC07F01F80FE03F80FE03F80FE03F80FE03F80FE03F80FE03F807F01FC07F01FC07F01FC03F80FE03F80FE01FC07F01FC03F80FE03";

cyclonev_ram_block ram_block1a60(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a60_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a60.clk0_core_clock_enable = "ena0";
defparam ram_block1a60.clk0_input_clock_enable = "ena0";
defparam ram_block1a60.clk0_output_clock_enable = "ena0";
defparam ram_block1a60.data_interleave_offset_in_bits = 1;
defparam ram_block1a60.data_interleave_width_in_bits = 1;
defparam ram_block1a60.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a60.init_file_layout = "port_a";
defparam ram_block1a60.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a60.operation_mode = "rom";
defparam ram_block1a60.port_a_address_clear = "none";
defparam ram_block1a60.port_a_address_width = 13;
defparam ram_block1a60.port_a_data_out_clear = "none";
defparam ram_block1a60.port_a_data_out_clock = "clock0";
defparam ram_block1a60.port_a_data_width = 1;
defparam ram_block1a60.port_a_first_address = 16384;
defparam ram_block1a60.port_a_first_bit_number = 12;
defparam ram_block1a60.port_a_last_address = 24575;
defparam ram_block1a60.port_a_logical_ram_depth = 65536;
defparam ram_block1a60.port_a_logical_ram_width = 24;
defparam ram_block1a60.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a60.ram_block_type = "auto";
defparam ram_block1a60.mem_init3 = "03F80FE03FC07F01FE03F80FF01FC03F80FE01FC07F80FE01FC07F80FE01FC03F80FF01FE03F807F00FE01FC03F80FF01FE03FC07F80FF01FE01FC03F807F00FF01FE03FC03F807F00FF01FE01FC03FC07F807F80FF00FE01FE01FC03FC03FC07F807F807F00FF00FF00FF01FE01FE01FE01FE01FE01FE01FC03FC03FC03FC03FE01FE01FE01FE01FE01FE01FE00FF00FF00FF007F807F807FC03FC03FE01FE01FF00FF007F807FC03FC01FE01FF00FF807F803FC01FE00FF007F803FC01FE00FF007F803FE01FF00FF803FC01FF00FF803FE01FF007F803FE00FF807FC01FF007FC03FE00FF803FE00FF803FE00FF803FE00FF803FE00FF803FE00FF801FF00";
defparam ram_block1a60.mem_init2 = "7FC01FF003FE00FF801FF007FC00FF803FF007FE00FF801FF003FE007FC00FF801FF003FE007FC00FFC01FF801FF003FF007FE007FE00FFC00FFC00FFC01FF801FF801FF801FF801FF801FF801FF801FF800FFC00FFC00FFC007FE007FF003FF003FF801FFC00FFC007FE003FF001FF800FFE007FF001FF800FFE007FF001FFC00FFE003FF800FFE003FF800FFE003FF800FFE003FF800FFF001FFC007FF800FFE001FFC007FF800FFF001FFE003FFC007FF8007FF000FFF000FFF001FFE001FFE001FFE001FFE001FFE001FFE000FFF000FFF0007FF8007FFC003FFE001FFF000FFF8003FFC001FFF000FFF8003FFE000FFF8003FFE000FFF8003FFF0007FFC";
defparam ram_block1a60.mem_init1 = "001FFF8003FFF0007FFE000FFFC000FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFF8000FFFC0007FFE0003FFF0001FFFC000FFFE0003FFF8000FFFE0003FFFC0007FFF0000FFFE0003FFFC0003FFF80007FFF80007FFF80007FFF80007FFFC0003FFFE0001FFFF0000FFFF80003FFFE0000FFFF80001FFFF00007FFFE0000FFFFC0000FFFFC0000FFFFC0000FFFFE00007FFFF00003FFFF80000FFFFE00003FFFFC00007FFFF80000FFFFF00000FFFFF000007FFFF800003FFFFC00001FFFFF800003FFFFE000007FFFFE000007FFFFE000007FFFFF000001FFFFFC000007FFFFF8000007FFFFF8000007FFFFFC000003FFFFFE0000007FFFFFE0000";
defparam ram_block1a60.mem_init0 = "007FFFFFE0000003FFFFFF8000000FFFFFFF00000007FFFFFF80000003FFFFFFF00000003FFFFFFF80000000FFFFFFFF00000000FFFFFFFF800000001FFFFFFFF8000000007FFFFFFFF8000000003FFFFFFFFF0000000001FFFFFFFFFE0000000000FFFFFFFFFFE00000000000FFFFFFFFFFFC000000000003FFFFFFFFFFFF00000000000007FFFFFFFFFFFFF8000000000000007FFFFFFFFFFFFFFF800000000000000001FFFFFFFFFFFFFFFFFFF0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a84(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a84_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a84.clk0_core_clock_enable = "ena0";
defparam ram_block1a84.clk0_input_clock_enable = "ena0";
defparam ram_block1a84.clk0_output_clock_enable = "ena0";
defparam ram_block1a84.data_interleave_offset_in_bits = 1;
defparam ram_block1a84.data_interleave_width_in_bits = 1;
defparam ram_block1a84.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a84.init_file_layout = "port_a";
defparam ram_block1a84.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a84.operation_mode = "rom";
defparam ram_block1a84.port_a_address_clear = "none";
defparam ram_block1a84.port_a_address_width = 13;
defparam ram_block1a84.port_a_data_out_clear = "none";
defparam ram_block1a84.port_a_data_out_clock = "clock0";
defparam ram_block1a84.port_a_data_width = 1;
defparam ram_block1a84.port_a_first_address = 24576;
defparam ram_block1a84.port_a_first_bit_number = 12;
defparam ram_block1a84.port_a_last_address = 32767;
defparam ram_block1a84.port_a_logical_ram_depth = 65536;
defparam ram_block1a84.port_a_logical_ram_width = 24;
defparam ram_block1a84.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a84.ram_block_type = "auto";
defparam ram_block1a84.mem_init3 = "07C1F07C1F07C0F83E0F83E0F83F07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F07E0F83E0F83E0FC1F07C1F07C1F03E0F83E0F83E07C1F07C1F07C0F83E0F83E0F83F07C1F07C1F07E0F83E0F83E07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F83E0F83E0F81F07C1F07C1F83E0F83E0F81F07C1F07C1F83E0F83E0F81F07C1F07C0F83E0F83E07C1F07C1F07E0F83E0F83F07C1F07C1F83E0F83E07C1F07C1F03E0F83E0FC1F07C1F07E0F83E0F81F07C1F07E0F83E0F81F07C1F07E0F83E0FC1F07C1F03E0F83E0FC1F07C1F83E0F83F07C1F07E0F83E0F81F07C1F03E0F83F07C1F07E0F83E0FC1F07C1F83E0F81F07C1F03E0F83F07C1F03E0F83E07";
defparam ram_block1a84.mem_init2 = "C1F07E0F83E07C1F07E0F83E07C1F07E0F83E07C1F03E0F83F07C1F03E0F81F07C1F83E0FC1F07C0F83E07C1F07E0F83F07C1F83E0FC1F07E0F83E07C1F03E0F81F07C0F83F07C1F83E0FC1F07E0F83F07C1F83E07C1F03E0F81F07E0F83F07C0F83E07C1F83E0FC1F03E0FC1F07E0F81F07E0F83F07C0F83F07C0F83F07C0F83E07C1F83E07C1F83E07C1F83E07C1F83E07C0F83F07C0F83F07C0F83F07E0F81F07E0F81F03E0FC1F03E07C1F83E07C0F83F07E0F81F03E0FC1F83E07C0F83F07E0F81F03E0FC1F83F07C0F81F03E0FC1F83F07E0F81F03E07C0F83F07E0FC1F83F07C0F81F03E07C0F81F03E07C0F83F07E0FC1F83F07E0FC1F83F07E0FC1F";
defparam ram_block1a84.mem_init1 = "83F03E07C0F81F03E07C0F81F03E07E0FC1F83F07E0FC0F81F03E07C0FC1F83F07E07C0F81F03F07E0FC0F81F03F07E0FC0F81F03F07E0FC0F81F83F07E07C0FC1F83F03E07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0F81F83F03F07E07C0FC1F81F83F03E07E07C0FC0F81F83F03F07E07E0FC0FC1F81F83F03F03E07E07C0FC0FC1F81F83F03F03E07E07E07C0FC0FC1F81F81F83F03F03F07E07E07E07C0FC0FC0FC1F81F81F81F83F03F03F03F03F07E07E07E07E07E07E0FC0FC0FC0FC0FC0FC0FC0FC0FC0F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81FC0FC0FC0FC0FC0FC0FC0FC0FC0FC07E07E07E07E07E07F03F03F03F03F01F";
defparam ram_block1a84.mem_init0 = "81F81F81F80FC0FC0FC07E07E07E03F03F03F01F81F81FC0FC0FC07E07E07F03F03F81F81FC0FC0FE07E07F03F03F81F80FC0FC07E07F03F01F81FC0FC07E07F03F01F81FC0FC07E07F03F81F80FC07E07F03F81F80FC07E03F03F81FC0FE07F03F01F80FC07E03F01F80FC07E03F01F80FC07F03F81FC0FE07F03F80FC07E03F81FC0FE03F01F80FE07F01F80FC07F03F80FC07F03F80FC07F01F80FE07F01FC0FE03F01FC07E03F80FE07F01FC0FE03F80FC07F01FC07E03F80FE03F01FC07F01FC07E03F80FE03F80FE03F80FE07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F80FE03F80FE03F80FE03FC07F01FC07F01FE03F80FE03FC07F01FC";

cyclonev_ram_block ram_block1a12(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "rom";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "clock0";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 8191;
defparam ram_block1a12.port_a_logical_ram_depth = 65536;
defparam ram_block1a12.port_a_logical_ram_width = 24;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init3 = "7F01FC07F80FE03F80FF01FC07F01FC07F80FE03F80FE03F80FE03FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC0FE03F80FE03F80FE03F80FC07F01FC07F01F80FE03F80FC07F01FC07E03F80FE07F01FC0FE03F80FC07F01F80FE07F01FC0FE03F01FC07E03F81FC07E03F81FC07E03F01FC0FE03F01F80FE07F03F80FC07E03F81FC0FE07F03F81FC07E03F01F80FC07E03F01F80FC07E03F01F81FC0FE07F03F81F80FC07E03F03F81FC0FC07E03F03F81FC0FC07E07F03F01F81FC0FC07E07F03F01F81FC0FC07E07E03F03F81F81FC0FC0FE07E07F03F03F81F81FC0FC0FC07E07E07F03F03F01F81F81F80FC0FC0FC07E07E07E03F03F03F03";
defparam ram_block1a12.mem_init2 = "F01F81F81F81F81FC0FC0FC0FC0FC0FC07E07E07E07E07E07E07E07E07E07F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03E07E07E07E07E07E07E07E07E07E0FC0FC0FC0FC0FC0FC1F81F81F81F81F83F03F03F03F07E07E07E07C0FC0FC0FC1F81F81F83F03F03F07E07E07C0FC0FC0F81F81F83F03F07E07E07C0FC0F81F81F83F03F07E07E0FC0FC1F81F83F03E07E07C0FC0F81F83F03F07E07C0FC1F81F83F03E07E0FC0F81F83F03E07E0FC0F81F83F03E07E0FC0F81F83F07E07C0FC1F83F03E07E0FC1F81F03E07E0FC1F81F03E07E0FC1F81F03E07C0FC1F83F07E07C0F81F03E07E0FC1F83F07E0FC0F81F03E07C0F81F03E07C0F81F83";
defparam ram_block1a12.mem_init1 = "F07E0FC1F83F07E0FC1F83F07E0FC1F83E07C0F81F03E07C0F81F03E07C1F83F07E0FC1F83E07C0F81F03E0FC1F83F07E0F81F03E07C1F83F07E0F81F03E0FC1F83E07C0F83F07E0F81F03E0FC1F83E07C0F83F07C0F81F07E0F81F03E0FC1F03E0FC1F83E07C1F83E07C1F83E07C0F83F07C0F83F07C0F83F07C0F83F07C0F83E07C1F83E07C1F83E07C1F83E0FC1F03E0FC1F07E0F81F07E0F83F07C0F83E07C1F83E0FC1F03E0F81F07C0F83F07C1F83E0FC1F07E0F83F07C1F83E07C1F03E0F81F07C0F83E0FC1F07E0F83F07C1F83E0FC1F07C0F83E07C1F07E0F83F07C1F03E0F81F07C1F83E0F81F07C0F83E0FC1F07C0F83E0FC1F07C0F83E0FC1F07";
defparam ram_block1a12.mem_init0 = "C0F83E0F81F07C1F83E0F81F07C1F03E0F83F07C1F07E0F83E0FC1F07C1F83E0F81F07C1F03E0F83E0FC1F07C1F83E0F83F07C1F07E0F83E0F81F07C1F07E0F83E0FC1F07C1F03E0F83E0FC1F07C1F03E0F83E0FC1F07C1F07E0F83E0F81F07C1F07C0F83E0F83F07C1F07C1F83E0F83E0FC1F07C1F07C0F83E0F83E07C1F07C1F03E0F83E0F83F07C1F07C1F03E0F83E0F83F07C1F07C1F03E0F83E0F83F07C1F07C1F03E0F83E0F83E07C1F07C1F07C0F83E0F83E0FC1F07C1F07C1F83E0F83E0F83E07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F07E0F83E0F83E0FC1F07C1F07C1F03E0F83E0F83E07C1F07C1F07C1F83E0F83E0F83E07C1F07C1F07C0";

cyclonev_ram_block ram_block1a36(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a36_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a36.clk0_core_clock_enable = "ena0";
defparam ram_block1a36.clk0_input_clock_enable = "ena0";
defparam ram_block1a36.clk0_output_clock_enable = "ena0";
defparam ram_block1a36.data_interleave_offset_in_bits = 1;
defparam ram_block1a36.data_interleave_width_in_bits = 1;
defparam ram_block1a36.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a36.init_file_layout = "port_a";
defparam ram_block1a36.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a36.operation_mode = "rom";
defparam ram_block1a36.port_a_address_clear = "none";
defparam ram_block1a36.port_a_address_width = 13;
defparam ram_block1a36.port_a_data_out_clear = "none";
defparam ram_block1a36.port_a_data_out_clock = "clock0";
defparam ram_block1a36.port_a_data_width = 1;
defparam ram_block1a36.port_a_first_address = 8192;
defparam ram_block1a36.port_a_first_bit_number = 12;
defparam ram_block1a36.port_a_last_address = 16383;
defparam ram_block1a36.port_a_logical_ram_depth = 65536;
defparam ram_block1a36.port_a_logical_ram_width = 24;
defparam ram_block1a36.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a36.ram_block_type = "auto";
defparam ram_block1a36.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000001FFFFFFFFFFFFFFFFFFF000000000000000003FFFFFFFFFFFFFFFC000000000000003FFFFFFFFFFFFFC0000000000001FFFFFFFFFFFF8000000000007FFFFFFFFFFE00000000000FFFFFFFFFFE0000000000FFFFFFFFFF0000000001FFFFFFFFF8000000003FFFFFFFFC000000003FFFFFFFF000000003FFFFFFFE00000001FFFFFFFE00000003FFFFFFF80000001FFFFFFF80000003FFFFFFC0000001FFFFFFE0000003FFFFFF8000000FFFFFFC00";
defparam ram_block1a36.mem_init2 = "0000FFFFFFC000000FFFFFF8000007FFFFFC000003FFFFFC000003FFFFFC000007FFFFF000001FFFFFC00000FFFFFC00000FFFFFC00000FFFFF800003FFFFF000007FFFF800003FFFFC00001FFFFE00001FFFFE00003FFFFC00007FFFF80000FFFFE00003FFFF80001FFFFC0000FFFFE00007FFFE00007FFFE00007FFFE0000FFFFC0001FFFF00003FFFE0000FFFF80003FFFE0001FFFF0000FFFF80007FFFC0003FFFC0003FFFC0003FFFC0003FFF80007FFF8000FFFE0001FFFC0007FFF8000FFFE0003FFF8000FFFE0007FFF0001FFF8000FFFC0007FFE0003FFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFE0007FFE000FFFC001FFF8003FFF000";
defparam ram_block1a36.mem_init1 = "7FFC001FFF8003FFE000FFF8003FFE000FFF8003FFE001FFF0007FF8003FFE001FFF000FFF8007FFC003FFC001FFE001FFE000FFF000FFF000FFF000FFF000FFF000FFF001FFE001FFE001FFC003FFC007FF800FFF001FFE003FFC007FF000FFE003FFC007FF001FFE003FF800FFE003FF800FFE003FF800FFE003FF800FFE007FF001FFC00FFE003FF001FFC00FFE003FF001FF800FFC007FE007FF003FF801FF801FFC00FFC007FE007FE007FE003FF003FF003FF003FF003FF003FF003FF003FF007FE007FE007FE00FFC00FFC01FF801FF003FF007FE007FC00FF801FF003FE007FC00FF801FF003FE00FFC01FF803FE007FC01FF003FE00FF801FF007FC";
defparam ram_block1a36.mem_init0 = "01FF003FE00FF803FE00FF803FE00FF803FE00FF803FE00FF803FE00FF807FC01FF007FC03FE00FF803FC01FF00FF803FE01FF007F803FE01FF00FF803FC01FE00FF007F803FC01FE00FF007F803FC03FE01FF00FF007F807FC03FC01FE01FF00FF00FF807F807FC03FC03FC01FE01FE01FE00FF00FF00FF00FF00FF00FF00FF807F807F807F807F00FF00FF00FF00FF00FF00FF01FE01FE01FE01FC03FC03FC07F807F807F00FF00FE01FE03FC03FC07F807F00FF01FE01FC03F807F80FF01FE01FC03F807F00FF01FE03FC07F80FF01FE03F807F00FE01FC03F80FF01FE03F807F00FE03FC07F00FE03FC07F00FE03F807F01FE03F80FF01FC07F80FE03F80";

cyclonev_ram_block ram_block1a109(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a109_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a109.clk0_core_clock_enable = "ena0";
defparam ram_block1a109.clk0_input_clock_enable = "ena0";
defparam ram_block1a109.clk0_output_clock_enable = "ena0";
defparam ram_block1a109.data_interleave_offset_in_bits = 1;
defparam ram_block1a109.data_interleave_width_in_bits = 1;
defparam ram_block1a109.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a109.init_file_layout = "port_a";
defparam ram_block1a109.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a109.operation_mode = "rom";
defparam ram_block1a109.port_a_address_clear = "none";
defparam ram_block1a109.port_a_address_width = 13;
defparam ram_block1a109.port_a_data_out_clear = "none";
defparam ram_block1a109.port_a_data_out_clock = "clock0";
defparam ram_block1a109.port_a_data_width = 1;
defparam ram_block1a109.port_a_first_address = 32768;
defparam ram_block1a109.port_a_first_bit_number = 13;
defparam ram_block1a109.port_a_last_address = 40959;
defparam ram_block1a109.port_a_logical_ram_depth = 65536;
defparam ram_block1a109.port_a_logical_ram_width = 24;
defparam ram_block1a109.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a109.ram_block_type = "auto";
defparam ram_block1a109.mem_init3 = "8001FFF8000FFFC000FFFE0007FFE0007FFF0003FFF0003FFF0003FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFF0003FFF0003FFF0003FFF0007FFE0007FFE000FFFC000FFF8001FFF8003FFF0007FFE000FFFC000FFF8001FFF0007FFE000FFFC001FFF8003FFE0007FFC001FFF8003FFE000FFFC001FFF0007FFC000FFF8003FFE000FFF8003FFE0007FFC001FFF0007FFC001FFF0007FFC001FFE000FFF8003FFE000FFF8003FFC001FFF0007FFC003FFE000FFF8007FFC001FFE000FFF8007FFC001FFE000FFF8007FFC003FFE001FFF000FFF8007FFC003FFE001FFF000FFF8007FF8003FFC001FFE001FFF000FFF0007FF8007FFC003FFC003";
defparam ram_block1a109.mem_init2 = "FFE001FFE001FFE000FFF000FFF000FFF8007FF8007FF8007FF8007FF8007FFC003FFC003FFC003FFC003FFC003FFC003FFC003FFC007FF8007FF8007FF8007FF8007FF000FFF000FFF000FFE001FFE001FFE003FFC003FFC007FF8007FF800FFF000FFE001FFE003FFC003FF8007FF800FFF000FFE001FFC003FF8007FF800FFF001FFE003FFC007FF800FFF001FFE003FFC007FF800FFF001FFC003FF8007FF001FFE003FFC007FF000FFE003FFC007FF000FFE003FFC007FF000FFE003FF8007FF001FFC003FF800FFE001FFC007FF001FFE003FF800FFE001FFC007FF001FFC007FF800FFE003FF800FFE003FF800FFF001FFC007FF001FFC007FF001FFC";
defparam ram_block1a109.mem_init1 = "007FF001FFC007FF001FFC007FF001FFC007FF001FFC007FF001FFC007FE003FF800FFE003FF800FFE003FF001FFC007FF001FFC007FE003FF800FFE003FF001FFC007FF003FF800FFE003FF001FFC007FF003FF800FFE007FF001FFC00FFE003FF001FFC007FE003FF801FFC007FF003FF800FFC007FF003FF800FFC007FF003FF801FFC007FE003FF801FFC00FFE003FF001FF800FFE007FF003FF800FFC007FE003FF001FFC00FFE007FF003FF801FFC00FFE007FF003FF801FFC007FE003FF001FF800FFC00FFE007FF003FF801FFC00FFE007FF003FF801FF800FFC007FE003FF001FF801FFC00FFE007FF003FF001FF800FFC00FFE007FF003FF001FF8";
defparam ram_block1a109.mem_init0 = "00FFC00FFE007FE003FF001FF801FFC00FFC007FE007FF003FF001FF801FFC00FFE007FE003FF003FF001FF801FFC00FFC007FE007FF003FF001FF801FF800FFC00FFE007FE003FF003FF001FF801FFC00FFC00FFE007FE007FF003FF001FF801FF800FFC00FFC007FE007FE003FF003FF001FF801FF800FFC00FFC007FE007FE003FF003FF003FF801FF801FFC00FFC00FFC007FE007FE003FF003FF003FF801FF801FFC00FFC00FFC007FE007FE007FF003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE007FF003FF003FF001FF801FF801FF800FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF801FFC00FFC00FFC007FE007FE007FE";

cyclonev_ram_block ram_block1a133(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a133_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a133.clk0_core_clock_enable = "ena0";
defparam ram_block1a133.clk0_input_clock_enable = "ena0";
defparam ram_block1a133.clk0_output_clock_enable = "ena0";
defparam ram_block1a133.data_interleave_offset_in_bits = 1;
defparam ram_block1a133.data_interleave_width_in_bits = 1;
defparam ram_block1a133.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a133.init_file_layout = "port_a";
defparam ram_block1a133.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a133.operation_mode = "rom";
defparam ram_block1a133.port_a_address_clear = "none";
defparam ram_block1a133.port_a_address_width = 13;
defparam ram_block1a133.port_a_data_out_clear = "none";
defparam ram_block1a133.port_a_data_out_clock = "clock0";
defparam ram_block1a133.port_a_data_width = 1;
defparam ram_block1a133.port_a_first_address = 40960;
defparam ram_block1a133.port_a_first_bit_number = 13;
defparam ram_block1a133.port_a_last_address = 49151;
defparam ram_block1a133.port_a_logical_ram_depth = 65536;
defparam ram_block1a133.port_a_logical_ram_width = 24;
defparam ram_block1a133.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a133.ram_block_type = "auto";
defparam ram_block1a133.mem_init3 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000FFFFFFFFFFFFFFFFFFFFF00000000000000000001FFFFFFFFFFFFFFFFFFC000000000000000003FFFFFFFFFFFFFFFFC0000000000000001FFFFFFFFFFFFFFFC000000000000001FFFFFFFFFFFFFFC00000000000001FFFFFFFFFFFFFC0000000000000FFFFFFFFF";
defparam ram_block1a133.mem_init2 = "FFFF0000000000000FFFFFFFFFFFF8000000000003FFFFFFFFFFFC000000000007FFFFFFFFFFE00000000000FFFFFFFFFFF00000000000FFFFFFFFFFC00000000007FFFFFFFFFC0000000001FFFFFFFFFE0000000003FFFFFFFFF8000000000FFFFFFFFFC000000001FFFFFFFFF0000000007FFFFFFFF8000000007FFFFFFFF000000001FFFFFFFFC00000000FFFFFFFFC00000001FFFFFFFF000000007FFFFFFFC00000003FFFFFFFC00000003FFFFFFF80000000FFFFFFFE00000007FFFFFFF00000003FFFFFFF00000007FFFFFFE0000000FFFFFFF80000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000003FFFFFF8000000FFFFFFE0000003FFFFFF";
defparam ram_block1a133.mem_init1 = "8000001FFFFFFC000000FFFFFFC000000FFFFFFC000001FFFFFF8000003FFFFFE000000FFFFFF8000003FFFFFE000001FFFFFF000000FFFFFF000000FFFFFF000000FFFFFE000001FFFFFE000003FFFFF800000FFFFFE000003FFFFF800000FFFFFC000007FFFFE000003FFFFF000003FFFFF000003FFFFF000003FFFFF000007FFFFE00000FFFFFC00001FFFFF000003FFFFE00000FFFFF800007FFFFC00001FFFFE00000FFFFF800007FFFF800003FFFFC00003FFFFC00003FFFFC00003FFFFC00007FFFF800007FFFF00000FFFFE00001FFFFC00007FFFF80000FFFFE00003FFFF80000FFFFE00003FFFF00001FFFFC00007FFFE00003FFFF00001FFFF800";
defparam ram_block1a133.mem_init0 = "01FFFFC0000FFFFC0000FFFFC0000FFFFC0000FFFFC0000FFFFC0000FFFF80001FFFF80003FFFF00003FFFE0000FFFFC0001FFFF80003FFFE0000FFFFC0001FFFF00007FFFC0001FFFF00007FFFC0003FFFE0000FFFF80007FFFC0001FFFE0000FFFF00007FFF80003FFFC0001FFFE0001FFFF0000FFFF0000FFFF0000FFFF00007FFF80007FFF8000FFFF0000FFFF0000FFFF0001FFFE0001FFFE0003FFFC0007FFF80007FFF0000FFFE0003FFFC0007FFF8000FFFE0001FFFC0007FFF0001FFFE0003FFF8000FFFE0003FFF8000FFFE0003FFF8000FFFE0003FFF0001FFFC0007FFF0003FFF8000FFFC0007FFF0003FFF8001FFFC000FFFE0007FFF0003FFF";

cyclonev_ram_block ram_block1a157(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a157_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a157.clk0_core_clock_enable = "ena0";
defparam ram_block1a157.clk0_input_clock_enable = "ena0";
defparam ram_block1a157.clk0_output_clock_enable = "ena0";
defparam ram_block1a157.data_interleave_offset_in_bits = 1;
defparam ram_block1a157.data_interleave_width_in_bits = 1;
defparam ram_block1a157.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a157.init_file_layout = "port_a";
defparam ram_block1a157.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a157.operation_mode = "rom";
defparam ram_block1a157.port_a_address_clear = "none";
defparam ram_block1a157.port_a_address_width = 13;
defparam ram_block1a157.port_a_data_out_clear = "none";
defparam ram_block1a157.port_a_data_out_clock = "clock0";
defparam ram_block1a157.port_a_data_width = 1;
defparam ram_block1a157.port_a_first_address = 49152;
defparam ram_block1a157.port_a_first_bit_number = 13;
defparam ram_block1a157.port_a_last_address = 57343;
defparam ram_block1a157.port_a_logical_ram_depth = 65536;
defparam ram_block1a157.port_a_logical_ram_width = 24;
defparam ram_block1a157.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a157.ram_block_type = "auto";
defparam ram_block1a157.mem_init3 = "FFF8001FFFC000FFFE0007FFF0003FFF8001FFFC0007FFE0003FFF8001FFFC0007FFF0001FFF8000FFFE0003FFF8000FFFE0003FFF8000FFFE0003FFF8000FFFF0001FFFC0007FFF0000FFFE0003FFFC0007FFF8000FFFE0001FFFC0003FFFC0007FFF8000FFFF0000FFFF0001FFFE0001FFFE0001FFFE0003FFFC0003FFFC0001FFFE0001FFFE0001FFFE0001FFFF0000FFFF00007FFF80003FFFC0001FFFE0000FFFF00007FFFC0003FFFE0000FFFF80007FFFC0001FFFF00007FFFC0001FFFF00007FFFE0000FFFF80003FFFF00007FFFE0000FFFF80001FFFF80003FFFF00003FFFE00007FFFE00007FFFE00007FFFE00007FFFE00007FFFE00007FFFF00";
defparam ram_block1a157.mem_init2 = "003FFFF00001FFFF80000FFFFC00007FFFF00001FFFF80000FFFFE00003FFFF80000FFFFE00003FFFFC00007FFFF00000FFFFE00001FFFFC00003FFFFC00007FFFF800007FFFF800007FFFF800007FFFF800003FFFFC00003FFFFE00000FFFFF000007FFFFC00003FFFFE00000FFFFF800001FFFFF000007FFFFE00000FFFFFC00001FFFFF800001FFFFF800001FFFFF800001FFFFF800000FFFFFC000007FFFFE000003FFFFF800000FFFFFE000003FFFFF800000FFFFFF000000FFFFFE000001FFFFFE000001FFFFFE000001FFFFFF000000FFFFFF8000003FFFFFE000000FFFFFF8000003FFFFFF0000007FFFFFE0000007FFFFFE0000007FFFFFF0000003";
defparam ram_block1a157.mem_init1 = "FFFFFF8000000FFFFFFE0000003FFFFFF80000007FFFFFF80000007FFFFFF80000007FFFFFF80000003FFFFFFE0000000FFFFFFFC0000001FFFFFFF80000001FFFFFFFC0000000FFFFFFFE00000003FFFFFFF800000007FFFFFFF800000007FFFFFFFC00000001FFFFFFFF000000007FFFFFFFE000000007FFFFFFFF000000001FFFFFFFFC000000003FFFFFFFFC000000001FFFFFFFFF0000000007FFFFFFFFE0000000003FFFFFFFFF8000000000FFFFFFFFFF00000000007FFFFFFFFFC00000000007FFFFFFFFFE00000000001FFFFFFFFFFE00000000000FFFFFFFFFFFC000000000007FFFFFFFFFFF8000000000003FFFFFFFFFFFE0000000000001FFFF";
defparam ram_block1a157.mem_init0 = "FFFFFFFFE00000000000007FFFFFFFFFFFFF000000000000007FFFFFFFFFFFFFF0000000000000007FFFFFFFFFFFFFFF00000000000000007FFFFFFFFFFFFFFFF8000000000000000007FFFFFFFFFFFFFFFFFF00000000000000000001FFFFFFFFFFFFFFFFFFFFE00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a181(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a181_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a181.clk0_core_clock_enable = "ena0";
defparam ram_block1a181.clk0_input_clock_enable = "ena0";
defparam ram_block1a181.clk0_output_clock_enable = "ena0";
defparam ram_block1a181.data_interleave_offset_in_bits = 1;
defparam ram_block1a181.data_interleave_width_in_bits = 1;
defparam ram_block1a181.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a181.init_file_layout = "port_a";
defparam ram_block1a181.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a181.operation_mode = "rom";
defparam ram_block1a181.port_a_address_clear = "none";
defparam ram_block1a181.port_a_address_width = 13;
defparam ram_block1a181.port_a_data_out_clear = "none";
defparam ram_block1a181.port_a_data_out_clock = "clock0";
defparam ram_block1a181.port_a_data_width = 1;
defparam ram_block1a181.port_a_first_address = 57344;
defparam ram_block1a181.port_a_first_bit_number = 13;
defparam ram_block1a181.port_a_last_address = 65535;
defparam ram_block1a181.port_a_logical_ram_depth = 65536;
defparam ram_block1a181.port_a_logical_ram_width = 24;
defparam ram_block1a181.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a181.ram_block_type = "auto";
defparam ram_block1a181.mem_init3 = "FFC00FFC00FFC007FE007FE007FF003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE003FF003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE007FF003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE007FF003FF003FF801FF801FF800FFC00FFC007FE007FE007FF003FF003FF801FF801FF800FFC00FFC007FE007FE003FF003FF001FF801FF800FFC00FFC007FE007FE003FF003FF001FF801FFC00FFC00FFE007FE007FF003FF001FF801FF800FFC00FFE007FE003FF003FF001FF801FFC00FFC007FE007FF003FF001FF801FF800FFC00FFE007FF003FF001FF801FFC00FFC007FE007FF003FF001FF800FFC00FFE007FE00";
defparam ram_block1a181.mem_init2 = "3FF001FF801FFC00FFE007FE003FF001FF801FFC00FFE007FF003FF001FF800FFC007FE003FF003FF801FFC00FFE007FF003FF801FFC00FFE007FE003FF001FF800FFC007FF003FF801FFC00FFE007FF003FF801FFC00FFE007FF001FF800FFC007FE003FF801FFC00FFE003FF001FF800FFE007FF003FF800FFC007FF003FF801FFC007FE003FF801FFC007FE003FF801FFC007FF003FF800FFC007FF001FF800FFE007FF001FFC00FFE003FF801FFC007FF001FF800FFE003FF801FFC007FF001FF800FFE003FF800FFC007FF001FFC007FF001FF800FFE003FF800FFE003FF800FFC007FF001FFC007FF001FFC007FF001FFC007FF001FFC007FF001FFC00";
defparam ram_block1a181.mem_init1 = "7FF001FFC007FF001FFC007FF001FFE003FF800FFE003FF800FFE003FFC007FF001FFC007FF000FFE003FF800FFF001FFC007FF000FFE003FF8007FF001FFC003FF800FFE001FFC007FF800FFE001FFC007FF800FFE001FFC007FF800FFF001FFC003FF8007FF001FFE003FFC007FF800FFF001FFE003FFC007FF800FFF001FFE003FFC003FF8007FF000FFE001FFE003FFC003FF8007FF800FFF000FFE001FFE003FFC003FFC007FF8007FF800FFF000FFF000FFE001FFE001FFE001FFC003FFC003FFC003FFC003FFC007FF8007FF8007FF8007FF8007FF8007FF8007FF8007FFC003FFC003FFC003FFC003FFC003FFE001FFE001FFE000FFF000FFF000FFF";
defparam ram_block1a181.mem_init0 = "8007FF8007FFC003FFC001FFE001FFF000FFF0007FF8003FFC003FFE001FFF000FFF8007FFC003FFE001FFF000FFF8007FFC003FFE000FFF0007FFC003FFE000FFF0007FFC003FFE000FFF8007FFC001FFF0007FF8003FFE000FFF8003FFE000FFF0007FFC001FFF0007FFC001FFF0007FFC000FFF8003FFE000FFF8003FFE0007FFC001FFF0007FFE000FFF8003FFF0007FFC000FFF8003FFF0007FFE000FFFC001FFF0003FFE0007FFE000FFFC001FFF8003FFF0003FFE0007FFE000FFFC000FFFC001FFF8001FFF8001FFF8001FFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFF8001FFF8001FFF8001FFFC000FFFC000FFFE0007FFE0003FFF0003";

cyclonev_ram_block ram_block1a61(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a61_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a61.clk0_core_clock_enable = "ena0";
defparam ram_block1a61.clk0_input_clock_enable = "ena0";
defparam ram_block1a61.clk0_output_clock_enable = "ena0";
defparam ram_block1a61.data_interleave_offset_in_bits = 1;
defparam ram_block1a61.data_interleave_width_in_bits = 1;
defparam ram_block1a61.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a61.init_file_layout = "port_a";
defparam ram_block1a61.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a61.operation_mode = "rom";
defparam ram_block1a61.port_a_address_clear = "none";
defparam ram_block1a61.port_a_address_width = 13;
defparam ram_block1a61.port_a_data_out_clear = "none";
defparam ram_block1a61.port_a_data_out_clock = "clock0";
defparam ram_block1a61.port_a_data_width = 1;
defparam ram_block1a61.port_a_first_address = 16384;
defparam ram_block1a61.port_a_first_bit_number = 13;
defparam ram_block1a61.port_a_last_address = 24575;
defparam ram_block1a61.port_a_logical_ram_depth = 65536;
defparam ram_block1a61.port_a_logical_ram_width = 24;
defparam ram_block1a61.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a61.ram_block_type = "auto";
defparam ram_block1a61.mem_init3 = "0007FFE0003FFF0001FFF8000FFFC0007FFE0003FFF8001FFFC0007FFE0003FFF8000FFFE0007FFF0001FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFF0000FFFE0003FFF8000FFFF0001FFFC0003FFF80007FFF0001FFFE0003FFFC0003FFF80007FFF0000FFFF0000FFFE0001FFFE0001FFFE0001FFFC0003FFFC0003FFFE0001FFFE0001FFFE0001FFFE0000FFFF0000FFFF80007FFFC0003FFFE0001FFFF0000FFFF80003FFFC0001FFFF00007FFF80003FFFE0000FFFF80003FFFE0000FFFF80001FFFF00007FFFC0000FFFF80001FFFF00007FFFE00007FFFC0000FFFFC0001FFFF80001FFFF80001FFFF80001FFFF80001FFFF80001FFFF80000FF";
defparam ram_block1a61.mem_init2 = "FFC0000FFFFE00007FFFF00003FFFF80000FFFFE00007FFFF00001FFFFC00007FFFF00001FFFFC00003FFFF80000FFFFF00001FFFFE00003FFFFC00003FFFF800007FFFF800007FFFF800007FFFF800007FFFFC00003FFFFC00001FFFFF00000FFFFF800003FFFFC00001FFFFF000007FFFFE00000FFFFF800001FFFFF000003FFFFE000007FFFFE000007FFFFE000007FFFFE000007FFFFF000003FFFFF800001FFFFFC000007FFFFF000001FFFFFC000007FFFFF000000FFFFFF000001FFFFFE000001FFFFFE000001FFFFFE000000FFFFFF0000007FFFFFC000001FFFFFF0000007FFFFFC000000FFFFFF8000001FFFFFF8000001FFFFFF8000000FFFFFFC";
defparam ram_block1a61.mem_init1 = "0000007FFFFFF0000001FFFFFFC0000007FFFFFF80000007FFFFFF80000007FFFFFF80000007FFFFFFC0000001FFFFFFF00000003FFFFFFE00000007FFFFFFE00000003FFFFFFF00000001FFFFFFFC00000007FFFFFFF800000007FFFFFFF800000003FFFFFFFE00000000FFFFFFFF800000001FFFFFFFF800000000FFFFFFFFE000000003FFFFFFFFC000000003FFFFFFFFE000000000FFFFFFFFF8000000001FFFFFFFFFC0000000007FFFFFFFFF0000000000FFFFFFFFFF80000000003FFFFFFFFFF80000000001FFFFFFFFFFE00000000001FFFFFFFFFFF000000000003FFFFFFFFFFF8000000000007FFFFFFFFFFFC000000000001FFFFFFFFFFFFE0000";
defparam ram_block1a61.mem_init0 = "000000001FFFFFFFFFFFFF80000000000000FFFFFFFFFFFFFF800000000000000FFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFF800000000000000007FFFFFFFFFFFFFFFFF8000000000000000000FFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a85(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a85_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a85.clk0_core_clock_enable = "ena0";
defparam ram_block1a85.clk0_input_clock_enable = "ena0";
defparam ram_block1a85.clk0_output_clock_enable = "ena0";
defparam ram_block1a85.data_interleave_offset_in_bits = 1;
defparam ram_block1a85.data_interleave_width_in_bits = 1;
defparam ram_block1a85.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a85.init_file_layout = "port_a";
defparam ram_block1a85.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a85.operation_mode = "rom";
defparam ram_block1a85.port_a_address_clear = "none";
defparam ram_block1a85.port_a_address_width = 13;
defparam ram_block1a85.port_a_data_out_clear = "none";
defparam ram_block1a85.port_a_data_out_clock = "clock0";
defparam ram_block1a85.port_a_data_width = 1;
defparam ram_block1a85.port_a_first_address = 24576;
defparam ram_block1a85.port_a_first_bit_number = 13;
defparam ram_block1a85.port_a_last_address = 32767;
defparam ram_block1a85.port_a_logical_ram_depth = 65536;
defparam ram_block1a85.port_a_logical_ram_width = 24;
defparam ram_block1a85.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a85.ram_block_type = "auto";
defparam ram_block1a85.mem_init3 = "003FF003FF003FF801FF801FF800FFC00FFC00FFC007FE007FE007FF003FF003FF001FF801FF801FFC00FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC007FE007FE007FF003FF003FF801FF801FF800FFC00FFC007FE007FE007FF003FF003FF801FF801FFC00FFC00FFE007FE007FF003FF003FF801FF801FFC00FFC00FFE007FE003FF003FF001FF801FF800FFC00FFE007FE007FF003FF001FF801FFC00FFC00FFE007FE003FF003FF801FF800FFC00FFE007FE007FF003FF001FF800FFC00FFE007FE003FF003FF801FF800FFC00FFE007FF003FF001FF801FF";
defparam ram_block1a85.mem_init2 = "C00FFE007FE003FF001FF801FFC00FFE007FE003FF001FF800FFC00FFE007FF003FF801FFC00FFC007FE003FF001FF800FFC007FE003FF001FF801FFC00FFE007FF003FF800FFC007FE003FF001FF800FFC007FE003FF001FF800FFE007FF003FF801FFC007FE003FF001FFC00FFE007FF001FF800FFC007FF003FF800FFC007FE003FF801FFC007FE003FF801FFC007FE003FF800FFC007FF003FF800FFE007FF001FF800FFE003FF001FFC007FE003FF800FFE007FF001FFC007FE003FF800FFE007FF001FFC007FF003FF800FFE003FF800FFE007FF001FFC007FF001FFC007FF003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF";
defparam ram_block1a85.mem_init1 = "800FFE003FF800FFE003FF800FFE001FFC007FF001FFC007FF001FFC003FF800FFE003FF800FFF001FFC007FF000FFE003FF800FFF001FFC007FF800FFE003FFC007FF001FFE003FF8007FF001FFE003FF8007FF001FFE003FF8007FF000FFE003FFC007FF800FFE001FFC003FF8007FF000FFE001FFC003FF8007FF000FFE001FFC003FFC007FF800FFF001FFE001FFC003FFC007FF8007FF000FFF001FFE001FFC003FFC003FF8007FF8007FF000FFF000FFF001FFE001FFE001FFE003FFC003FFC003FFC003FFC003FF8007FF8007FF8007FF8007FF8007FF8007FF8007FF8003FFC003FFC003FFC003FFC003FFC001FFE001FFE001FFF000FFF000FFF000";
defparam ram_block1a85.mem_init0 = "7FF8007FF8003FFC003FFE001FFE000FFF000FFF8007FFC003FFC001FFE000FFF0007FF8003FFC001FFE000FFF0007FF8003FFC001FFF000FFF8003FFC001FFF000FFF8003FFC001FFF0007FF8003FFE000FFF8007FFC001FFF0007FFC001FFF000FFF8003FFE000FFF8003FFE000FFF8003FFF0007FFC001FFF0007FFC001FFF8003FFE000FFF8001FFF0007FFC000FFF8003FFF0007FFC000FFF8001FFF0003FFE000FFFC001FFF8001FFF0003FFE0007FFC000FFFC001FFF8001FFF0003FFF0003FFE0007FFE0007FFE0007FFE000FFFC000FFFC000FFFC000FFFC000FFFC000FFFC0007FFE0007FFE0007FFE0003FFF0003FFF0001FFF8001FFFC000FFFC";

cyclonev_ram_block ram_block1a13(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "rom";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "clock0";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 8191;
defparam ram_block1a13.port_a_logical_ram_depth = 65536;
defparam ram_block1a13.port_a_logical_ram_width = 24;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init3 = "7FFE0007FFF0003FFF0001FFF8001FFF8000FFFC000FFFC000FFFC0007FFE0007FFE0007FFE0007FFE0007FFE0007FFE000FFFC000FFFC000FFFC000FFF8001FFF8001FFF0003FFF0007FFE0007FFC000FFF8001FFF0003FFF0007FFE000FFF8001FFF0003FFE0007FFC001FFF8003FFE0007FFC001FFF0003FFE000FFF8003FFF0007FFC001FFF0007FFC001FFF8003FFE000FFF8003FFE000FFF8003FFE001FFF0007FFC001FFF0007FFC003FFE000FFF8003FFC001FFF0007FF8003FFE001FFF0007FF8003FFE001FFF0007FF8003FFC001FFE000FFF0007FF8003FFC001FFE000FFF0007FF8007FFC003FFE001FFE000FFF000FFF8007FF8003FFC003FFC";
defparam ram_block1a13.mem_init2 = "001FFE001FFE001FFF000FFF000FFF0007FF8007FF8007FF8007FF8007FF8003FFC003FFC003FFC003FFC003FFC003FFC003FFC003FF8007FF8007FF8007FF8007FF800FFF000FFF000FFF001FFE001FFE001FFC003FFC003FF8007FF8007FF000FFF001FFE001FFC003FFC007FF8007FF000FFF001FFE003FFC007FF8007FF000FFE001FFC003FF8007FF000FFE001FFC003FF8007FF000FFE003FFC007FF800FFE001FFC003FF800FFF001FFC003FF800FFF001FFC003FF800FFF001FFC007FF800FFE003FFC007FF001FFE003FF800FFE001FFC007FF001FFE003FF800FFE003FF8007FF001FFC007FF001FFC007FF000FFE003FF800FFE003FF800FFE003";
defparam ram_block1a13.mem_init1 = "FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF801FFC007FF001FFC007FF001FFC00FFE003FF800FFE003FF801FFC007FF001FFC00FFE003FF800FFC007FF001FFC00FFE003FF800FFC007FF001FF800FFE003FF001FFC00FFE003FF801FFC007FE003FF800FFC007FF003FF800FFC007FF003FF800FFC007FE003FF801FFC007FE003FF001FFC00FFE007FF001FF800FFC007FF003FF801FFC00FFE003FF001FF800FFC007FE003FF001FF800FFC007FE003FF801FFC00FFE007FF003FF001FF800FFC007FE003FF001FF800FFC007FE007FF003FF801FFC00FFE007FE003FF001FF800FFC00FFE007FF003FF001FF800FFC00FFE007";
defparam ram_block1a13.mem_init0 = "FF003FF001FF801FFC00FFE007FE003FF003FF801FF800FFC00FFE007FE003FF001FF801FFC00FFC00FFE007FE003FF003FF801FF800FFC00FFE007FE007FF003FF001FF801FFC00FFC00FFE007FE003FF003FF001FF801FF800FFC00FFE007FE007FF003FF003FF801FF801FFC00FFC00FFE007FE007FF003FF003FF801FF801FFC00FFC00FFC007FE007FE003FF003FF003FF801FF801FFC00FFC00FFC007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE007FF003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE007FE003FF003FF003FF801FF801FF800";

cyclonev_ram_block ram_block1a37(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a37_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a37.clk0_core_clock_enable = "ena0";
defparam ram_block1a37.clk0_input_clock_enable = "ena0";
defparam ram_block1a37.clk0_output_clock_enable = "ena0";
defparam ram_block1a37.data_interleave_offset_in_bits = 1;
defparam ram_block1a37.data_interleave_width_in_bits = 1;
defparam ram_block1a37.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a37.init_file_layout = "port_a";
defparam ram_block1a37.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a37.operation_mode = "rom";
defparam ram_block1a37.port_a_address_clear = "none";
defparam ram_block1a37.port_a_address_width = 13;
defparam ram_block1a37.port_a_data_out_clear = "none";
defparam ram_block1a37.port_a_data_out_clock = "clock0";
defparam ram_block1a37.port_a_data_width = 1;
defparam ram_block1a37.port_a_first_address = 8192;
defparam ram_block1a37.port_a_first_bit_number = 13;
defparam ram_block1a37.port_a_last_address = 16383;
defparam ram_block1a37.port_a_logical_ram_depth = 65536;
defparam ram_block1a37.port_a_logical_ram_width = 24;
defparam ram_block1a37.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a37.ram_block_type = "auto";
defparam ram_block1a37.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFE0000000000000000003FFFFFFFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFE0000000000000003FFFFFFFFFFFFFFE000000000000003FFFFFFFFFFFFFE00000000000003FFFFFFFFFFFFF000000000";
defparam ram_block1a37.mem_init2 = "0000FFFFFFFFFFFFF0000000000007FFFFFFFFFFFC000000000003FFFFFFFFFFF800000000001FFFFFFFFFFF00000000000FFFFFFFFFFF00000000003FFFFFFFFFF80000000003FFFFFFFFFE0000000001FFFFFFFFFC0000000007FFFFFFFFF0000000003FFFFFFFFE000000000FFFFFFFFF8000000007FFFFFFFF800000000FFFFFFFFE000000003FFFFFFFF000000003FFFFFFFE00000000FFFFFFFF800000003FFFFFFFC00000003FFFFFFFC00000007FFFFFFF00000001FFFFFFF80000000FFFFFFFC0000000FFFFFFF80000001FFFFFFF00000007FFFFFFC0000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000007FFFFFF0000001FFFFFFC000000";
defparam ram_block1a37.mem_init1 = "7FFFFFE0000003FFFFFF0000003FFFFFF0000003FFFFFE0000007FFFFFC000001FFFFFF0000007FFFFFC000001FFFFFE000000FFFFFF000000FFFFFF000000FFFFFF000001FFFFFE000001FFFFFC000007FFFFF000001FFFFFC000007FFFFF000003FFFFF800001FFFFFC00000FFFFFC00000FFFFFC00000FFFFFC00000FFFFF800001FFFFF000003FFFFE00000FFFFFC00001FFFFF000007FFFF800003FFFFE00001FFFFF000007FFFF800007FFFFC00003FFFFC00003FFFFC00003FFFFC00003FFFF800007FFFF80000FFFFF00001FFFFE00003FFFF800007FFFF00001FFFFC00007FFFF00001FFFFC0000FFFFE00003FFFF80001FFFFC0000FFFFE00007FF";
defparam ram_block1a37.mem_init0 = "FE00003FFFF00003FFFF00003FFFF00003FFFF00003FFFF00003FFFF00007FFFE00007FFFC0000FFFFC0001FFFF00003FFFE00007FFFC0001FFFF00003FFFE0000FFFF80003FFFE0000FFFF80003FFFC0001FFFF00007FFF80003FFFE0001FFFF0000FFFF80007FFFC0003FFFE0001FFFE0000FFFF0000FFFF0000FFFF0000FFFF80007FFF80007FFF0000FFFF0000FFFF0000FFFE0001FFFE0001FFFC0003FFF80007FFF8000FFFF0001FFFC0003FFF80007FFF0001FFFE0003FFF8000FFFE0001FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFF0001FFFC000FFFE0003FFF8000FFFC0007FFF0003FFF8000FFFC0007FFE0003FFF0001FFF8000FFFC000";

cyclonev_ram_block ram_block1a110(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a110_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a110.clk0_core_clock_enable = "ena0";
defparam ram_block1a110.clk0_input_clock_enable = "ena0";
defparam ram_block1a110.clk0_output_clock_enable = "ena0";
defparam ram_block1a110.data_interleave_offset_in_bits = 1;
defparam ram_block1a110.data_interleave_width_in_bits = 1;
defparam ram_block1a110.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a110.init_file_layout = "port_a";
defparam ram_block1a110.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a110.operation_mode = "rom";
defparam ram_block1a110.port_a_address_clear = "none";
defparam ram_block1a110.port_a_address_width = 13;
defparam ram_block1a110.port_a_data_out_clear = "none";
defparam ram_block1a110.port_a_data_out_clock = "clock0";
defparam ram_block1a110.port_a_data_width = 1;
defparam ram_block1a110.port_a_first_address = 32768;
defparam ram_block1a110.port_a_first_bit_number = 14;
defparam ram_block1a110.port_a_last_address = 40959;
defparam ram_block1a110.port_a_logical_ram_depth = 65536;
defparam ram_block1a110.port_a_logical_ram_width = 24;
defparam ram_block1a110.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a110.ram_block_type = "auto";
defparam ram_block1a110.mem_init3 = "80000007FFFFFFC0000001FFFFFFE0000000FFFFFFF0000000FFFFFFF80000007FFFFFF80000007FFFFFF80000007FFFFFF0000000FFFFFFF0000000FFFFFFE0000001FFFFFFC0000007FFFFFF8000000FFFFFFE0000003FFFFFF8000000FFFFFFE0000003FFFFFF8000001FFFFFFC0000007FFFFFE0000003FFFFFF0000003FFFFFF8000001FFFFFF8000001FFFFFFC000000FFFFFFC000000FFFFFFC000001FFFFFF8000001FFFFFF8000003FFFFFF0000003FFFFFE0000007FFFFFC000001FFFFFF8000003FFFFFE0000007FFFFFC000001FFFFFF0000007FFFFFC000001FFFFFF0000007FFFFF8000003FFFFFE000000FFFFFF0000007FFFFFC000003FFF";
defparam ram_block1a110.mem_init2 = "FFE000001FFFFFE000000FFFFFF0000007FFFFF8000007FFFFF8000007FFFFFC000003FFFFFC000003FFFFFC000003FFFFFC000003FFFFF8000007FFFFF8000007FFFFF000000FFFFFF000001FFFFFE000001FFFFFC000003FFFFF8000007FFFFF000001FFFFFE000003FFFFF8000007FFFFF000001FFFFFC000007FFFFF800000FFFFFE000003FFFFF800000FFFFFE000003FFFFF800000FFFFFC000007FFFFF000001FFFFFC00000FFFFFE000003FFFFF000001FFFFFC00000FFFFFE000007FFFFF000003FFFFF800001FFFFFC00000FFFFFE000007FFFFE000003FFFFF000003FFFFF800001FFFFF800001FFFFF800000FFFFFC00000FFFFFC00000FFFFFC";
defparam ram_block1a110.mem_init1 = "00000FFFFFC00000FFFFFC00000FFFFFC00000FFFFFC00000FFFFFC00001FFFFF800001FFFFF800001FFFFF000003FFFFF000003FFFFE000007FFFFE00000FFFFFC00000FFFFF800001FFFFF000003FFFFF000007FFFFE00000FFFFFC00001FFFFF000003FFFFE000007FFFFC00000FFFFF800003FFFFF000007FFFFC00000FFFFF800003FFFFE000007FFFFC00001FFFFF000007FFFFE00000FFFFF800003FFFFE00000FFFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF000007FFFFC00001FFFFF00000FFFFF8";
defparam ram_block1a110.mem_init0 = "00003FFFFE00001FFFFF000007FFFFC00003FFFFE00000FFFFF000007FFFFC00001FFFFE00000FFFFF000007FFFFC00003FFFFE00000FFFFF000007FFFF800003FFFFE00001FFFFF00000FFFFF800003FFFFC00001FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF000007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFC00001FFFFE00000FFFFF00000FFFFF800007FFFFC00003FFFFC00001FFFFE00000FFFFF00000FFFFF800007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00003FFFFE00001FFFFE";

cyclonev_ram_block ram_block1a134(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a134_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a134.clk0_core_clock_enable = "ena0";
defparam ram_block1a134.clk0_input_clock_enable = "ena0";
defparam ram_block1a134.clk0_output_clock_enable = "ena0";
defparam ram_block1a134.data_interleave_offset_in_bits = 1;
defparam ram_block1a134.data_interleave_width_in_bits = 1;
defparam ram_block1a134.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a134.init_file_layout = "port_a";
defparam ram_block1a134.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a134.operation_mode = "rom";
defparam ram_block1a134.port_a_address_clear = "none";
defparam ram_block1a134.port_a_address_width = 13;
defparam ram_block1a134.port_a_data_out_clear = "none";
defparam ram_block1a134.port_a_data_out_clock = "clock0";
defparam ram_block1a134.port_a_data_width = 1;
defparam ram_block1a134.port_a_first_address = 40960;
defparam ram_block1a134.port_a_first_bit_number = 14;
defparam ram_block1a134.port_a_last_address = 49151;
defparam ram_block1a134.port_a_logical_ram_depth = 65536;
defparam ram_block1a134.port_a_logical_ram_width = 24;
defparam ram_block1a134.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a134.ram_block_type = "auto";
defparam ram_block1a134.mem_init3 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a134.mem_init2 = "FFFF00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000001FFFFFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFF80000000000000000003FFFFFFFFFFFFFFFFFF0000000000000000007FFFFFFFFFFFFFFFFF000000000000000003FFFFFFFFFFFFFFFFC0000000000000000FFFFFFFFFFFFFFFFC0000000000000003FFFFFFFFFFFFFFF8000000000000001FFFFFFFFFFFFFFF000000000000000FFFFFFFFFFFFFFE000000000000007FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFC00000000000007FFFFFFFFFFFFE0000000000000";
defparam ram_block1a134.mem_init1 = "7FFFFFFFFFFFFC0000000000003FFFFFFFFFFFFC0000000000007FFFFFFFFFFFE0000000000007FFFFFFFFFFFE000000000000FFFFFFFFFFFF000000000000FFFFFFFFFFFE000000000001FFFFFFFFFFF800000000001FFFFFFFFFFF800000000003FFFFFFFFFFE00000000000FFFFFFFFFFF00000000000FFFFFFFFFFF00000000001FFFFFFFFFFC0000000000FFFFFFFFFFE00000000007FFFFFFFFFC0000000001FFFFFFFFFF80000000007FFFFFFFFFC0000000003FFFFFFFFFC0000000003FFFFFFFFF8000000000FFFFFFFFFE0000000003FFFFFFFFF8000000001FFFFFFFFF8000000001FFFFFFFFF0000000003FFFFFFFFE000000000FFFFFFFFF800";
defparam ram_block1a134.mem_init0 = "0000003FFFFFFFFC000000003FFFFFFFFC000000003FFFFFFFFC000000007FFFFFFFF800000000FFFFFFFFE000000003FFFFFFFF800000001FFFFFFFFC00000000FFFFFFFFC00000000FFFFFFFFC00000001FFFFFFFF800000003FFFFFFFE00000000FFFFFFFF800000003FFFFFFFE00000000FFFFFFFF00000000FFFFFFFF000000007FFFFFFF80000000FFFFFFFF00000000FFFFFFFE00000001FFFFFFFC00000007FFFFFFF00000001FFFFFFFC00000007FFFFFFE00000003FFFFFFF00000001FFFFFFF80000001FFFFFFF80000001FFFFFFF80000001FFFFFFF00000003FFFFFFF00000007FFFFFFC0000000FFFFFFF80000003FFFFFFE0000000FFFFFFF";

cyclonev_ram_block ram_block1a158(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a158_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a158.clk0_core_clock_enable = "ena0";
defparam ram_block1a158.clk0_input_clock_enable = "ena0";
defparam ram_block1a158.clk0_output_clock_enable = "ena0";
defparam ram_block1a158.data_interleave_offset_in_bits = 1;
defparam ram_block1a158.data_interleave_width_in_bits = 1;
defparam ram_block1a158.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a158.init_file_layout = "port_a";
defparam ram_block1a158.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a158.operation_mode = "rom";
defparam ram_block1a158.port_a_address_clear = "none";
defparam ram_block1a158.port_a_address_width = 13;
defparam ram_block1a158.port_a_data_out_clear = "none";
defparam ram_block1a158.port_a_data_out_clock = "clock0";
defparam ram_block1a158.port_a_data_width = 1;
defparam ram_block1a158.port_a_first_address = 49152;
defparam ram_block1a158.port_a_first_bit_number = 14;
defparam ram_block1a158.port_a_last_address = 57343;
defparam ram_block1a158.port_a_logical_ram_depth = 65536;
defparam ram_block1a158.port_a_logical_ram_width = 24;
defparam ram_block1a158.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a158.ram_block_type = "auto";
defparam ram_block1a158.mem_init3 = "FFFFFFE0000000FFFFFFF80000003FFFFFFE00000007FFFFFFC0000001FFFFFFF80000001FFFFFFF00000003FFFFFFF00000003FFFFFFF00000003FFFFFFF00000001FFFFFFF80000000FFFFFFFC00000007FFFFFFF00000001FFFFFFFC00000007FFFFFFF00000000FFFFFFFE00000001FFFFFFFE00000003FFFFFFFC00000001FFFFFFFE00000001FFFFFFFE00000000FFFFFFFF800000003FFFFFFFE00000000FFFFFFFF800000003FFFFFFFF000000007FFFFFFFE000000007FFFFFFFE000000007FFFFFFFF000000003FFFFFFFF800000000FFFFFFFFE000000003FFFFFFFFC000000007FFFFFFFF8000000007FFFFFFFF8000000007FFFFFFFF8000000";
defparam ram_block1a158.mem_init2 = "003FFFFFFFFE000000000FFFFFFFFF8000000001FFFFFFFFF0000000003FFFFFFFFF0000000003FFFFFFFFF8000000000FFFFFFFFFE0000000003FFFFFFFFF80000000007FFFFFFFFF80000000007FFFFFFFFFC0000000003FFFFFFFFFF00000000007FFFFFFFFFC0000000000FFFFFFFFFFE00000000007FFFFFFFFFF00000000001FFFFFFFFFFE00000000001FFFFFFFFFFE00000000000FFFFFFFFFFF800000000003FFFFFFFFFFF000000000003FFFFFFFFFFF000000000000FFFFFFFFFFFE000000000001FFFFFFFFFFFE000000000000FFFFFFFFFFFFC000000000000FFFFFFFFFFFFC0000000000007FFFFFFFFFFFF80000000000007FFFFFFFFFFFFC";
defparam ram_block1a158.mem_init1 = "0000000000000FFFFFFFFFFFFFC00000000000007FFFFFFFFFFFFF800000000000007FFFFFFFFFFFFFC00000000000000FFFFFFFFFFFFFFE000000000000001FFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFF80000000000000007FFFFFFFFFFFFFFFE00000000000000007FFFFFFFFFFFFFFFF800000000000000001FFFFFFFFFFFFFFFFFC000000000000000001FFFFFFFFFFFFFFFFFF80000000000000000003FFFFFFFFFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFFFFF8000000000000000000001FFFFFFFFFFFFFFFFFFFFFF000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000001FFFF";
defparam ram_block1a158.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a182(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a182_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a182.clk0_core_clock_enable = "ena0";
defparam ram_block1a182.clk0_input_clock_enable = "ena0";
defparam ram_block1a182.clk0_output_clock_enable = "ena0";
defparam ram_block1a182.data_interleave_offset_in_bits = 1;
defparam ram_block1a182.data_interleave_width_in_bits = 1;
defparam ram_block1a182.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a182.init_file_layout = "port_a";
defparam ram_block1a182.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a182.operation_mode = "rom";
defparam ram_block1a182.port_a_address_clear = "none";
defparam ram_block1a182.port_a_address_width = 13;
defparam ram_block1a182.port_a_data_out_clear = "none";
defparam ram_block1a182.port_a_data_out_clock = "clock0";
defparam ram_block1a182.port_a_data_width = 1;
defparam ram_block1a182.port_a_first_address = 57344;
defparam ram_block1a182.port_a_first_bit_number = 14;
defparam ram_block1a182.port_a_last_address = 65535;
defparam ram_block1a182.port_a_logical_ram_depth = 65536;
defparam ram_block1a182.port_a_logical_ram_width = 24;
defparam ram_block1a182.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a182.ram_block_type = "auto";
defparam ram_block1a182.mem_init3 = "FFFFF00000FFFFF800007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC00003FFFFE00001FFFFE00000FFFFF000007FFFF800007FFFFC00003FFFFE00001FFFFE00000FFFFF000007FFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00001FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF000007FFFF800003FFFFE00001FFFFF00000FFFFF800003FFFFC00001FFFFE00000FFFFF800007FFFFC00001FFFFE00000FFFFF000007FFFFC00001FFFFE00000FFFFF800007FFFFC00001FFFFF00000FFFFF80000";
defparam ram_block1a182.mem_init2 = "3FFFFE00001FFFFF000007FFFFC00001FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFE00000FFFFF800003FFFFE00000FFFFFC00001FFFFF000007FFFFC00000FFFFF800003FFFFE000007FFFFC00001FFFFF800003FFFFE000007FFFFC00000FFFFF800001FFFFF000007FFFFE00000FFFFFC00001FFFFF800001FFFFF000003FFFFE000007FFFFE00000FFFFFC00000FFFFF800001FFFFF800001FFFFF000003FFFFF000003FFFFF000007FFFFE000007FFFFE000007FFFFE000007FFFFE000007FFFFE00000";
defparam ram_block1a182.mem_init1 = "7FFFFE000007FFFFE000007FFFFE000003FFFFF000003FFFFF000003FFFFF800001FFFFF800000FFFFFC00000FFFFFE000007FFFFF000003FFFFF800001FFFFFC00000FFFFFE000007FFFFF000001FFFFF800000FFFFFE000007FFFFF000001FFFFFC000007FFFFE000003FFFFF800000FFFFFE000003FFFFF800000FFFFFE000003FFFFFC000007FFFFF000001FFFFFC000003FFFFF800000FFFFFF000001FFFFFC000003FFFFF8000007FFFFF000000FFFFFF000001FFFFFE000001FFFFFC000003FFFFFC000003FFFFF8000007FFFFF8000007FFFFF8000007FFFFF8000007FFFFFC000003FFFFFC000003FFFFFC000001FFFFFE000000FFFFFF000000FFF";
defparam ram_block1a182.mem_init0 = "FFF8000007FFFFFC000001FFFFFE000000FFFFFF8000003FFFFFC000001FFFFFF0000007FFFFFC000001FFFFFF0000007FFFFFC000000FFFFFF8000003FFFFFF0000007FFFFFC000000FFFFFF8000001FFFFFF8000003FFFFFF0000003FFFFFF0000007FFFFFE0000007FFFFFE0000007FFFFFF0000003FFFFFF0000003FFFFFF8000001FFFFFF8000000FFFFFFC0000007FFFFFF0000003FFFFFF8000000FFFFFFE0000003FFFFFF8000000FFFFFFE0000003FFFFFFC0000007FFFFFF0000000FFFFFFE0000001FFFFFFE0000001FFFFFFC0000003FFFFFFC0000003FFFFFFC0000003FFFFFFE0000001FFFFFFE0000000FFFFFFF00000007FFFFFFC0000003";

cyclonev_ram_block ram_block1a62(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a62_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a62.clk0_core_clock_enable = "ena0";
defparam ram_block1a62.clk0_input_clock_enable = "ena0";
defparam ram_block1a62.clk0_output_clock_enable = "ena0";
defparam ram_block1a62.data_interleave_offset_in_bits = 1;
defparam ram_block1a62.data_interleave_width_in_bits = 1;
defparam ram_block1a62.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a62.init_file_layout = "port_a";
defparam ram_block1a62.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a62.operation_mode = "rom";
defparam ram_block1a62.port_a_address_clear = "none";
defparam ram_block1a62.port_a_address_width = 13;
defparam ram_block1a62.port_a_data_out_clear = "none";
defparam ram_block1a62.port_a_data_out_clock = "clock0";
defparam ram_block1a62.port_a_data_width = 1;
defparam ram_block1a62.port_a_first_address = 16384;
defparam ram_block1a62.port_a_first_bit_number = 14;
defparam ram_block1a62.port_a_last_address = 24575;
defparam ram_block1a62.port_a_logical_ram_depth = 65536;
defparam ram_block1a62.port_a_logical_ram_width = 24;
defparam ram_block1a62.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a62.ram_block_type = "auto";
defparam ram_block1a62.mem_init3 = "0000001FFFFFFF00000007FFFFFFC0000001FFFFFFF80000003FFFFFFE00000007FFFFFFE0000000FFFFFFFC0000000FFFFFFFC0000000FFFFFFFC0000000FFFFFFFE00000007FFFFFFF00000003FFFFFFF80000000FFFFFFFE00000003FFFFFFF80000000FFFFFFFF00000001FFFFFFFE00000001FFFFFFFC00000003FFFFFFFE00000001FFFFFFFE00000001FFFFFFFF000000007FFFFFFFC00000001FFFFFFFF000000007FFFFFFFC00000000FFFFFFFF800000001FFFFFFFF800000001FFFFFFFF800000000FFFFFFFFC000000007FFFFFFFF000000001FFFFFFFFC000000003FFFFFFFF8000000007FFFFFFFF8000000007FFFFFFFF8000000007FFFFFF";
defparam ram_block1a62.mem_init2 = "FFC000000001FFFFFFFFF0000000007FFFFFFFFE000000000FFFFFFFFFC000000000FFFFFFFFFC0000000007FFFFFFFFF0000000001FFFFFFFFFC0000000007FFFFFFFFF80000000007FFFFFFFFF80000000003FFFFFFFFFC0000000000FFFFFFFFFF80000000003FFFFFFFFFF00000000001FFFFFFFFFF80000000000FFFFFFFFFFE00000000001FFFFFFFFFFE00000000001FFFFFFFFFFF000000000007FFFFFFFFFFC00000000000FFFFFFFFFFFC00000000000FFFFFFFFFFFF000000000001FFFFFFFFFFFE000000000001FFFFFFFFFFFF0000000000003FFFFFFFFFFFF0000000000003FFFFFFFFFFFF80000000000007FFFFFFFFFFFF80000000000003";
defparam ram_block1a62.mem_init1 = "FFFFFFFFFFFFF00000000000003FFFFFFFFFFFFF800000000000007FFFFFFFFFFFFF800000000000003FFFFFFFFFFFFFF000000000000001FFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFFC0000000000000007FFFFFFFFFFFFFFF80000000000000001FFFFFFFFFFFFFFFF800000000000000007FFFFFFFFFFFFFFFFE000000000000000003FFFFFFFFFFFFFFFFFE0000000000000000007FFFFFFFFFFFFFFFFFFC0000000000000000000FFFFFFFFFFFFFFFFFFFF8000000000000000000007FFFFFFFFFFFFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFE0000";
defparam ram_block1a62.mem_init0 = "00000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a86(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a86_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a86.clk0_core_clock_enable = "ena0";
defparam ram_block1a86.clk0_input_clock_enable = "ena0";
defparam ram_block1a86.clk0_output_clock_enable = "ena0";
defparam ram_block1a86.data_interleave_offset_in_bits = 1;
defparam ram_block1a86.data_interleave_width_in_bits = 1;
defparam ram_block1a86.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a86.init_file_layout = "port_a";
defparam ram_block1a86.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a86.operation_mode = "rom";
defparam ram_block1a86.port_a_address_clear = "none";
defparam ram_block1a86.port_a_address_width = 13;
defparam ram_block1a86.port_a_data_out_clear = "none";
defparam ram_block1a86.port_a_data_out_clock = "clock0";
defparam ram_block1a86.port_a_data_width = 1;
defparam ram_block1a86.port_a_first_address = 24576;
defparam ram_block1a86.port_a_first_bit_number = 14;
defparam ram_block1a86.port_a_last_address = 32767;
defparam ram_block1a86.port_a_logical_ram_depth = 65536;
defparam ram_block1a86.port_a_logical_ram_width = 24;
defparam ram_block1a86.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a86.ram_block_type = "auto";
defparam ram_block1a86.mem_init3 = "00000FFFFF000007FFFF800007FFFFC00003FFFFC00001FFFFE00000FFFFF00000FFFFF800007FFFFC00003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00001FFFFE00000FFFFF000007FFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00001FFFFE00000FFFFF000007FFFFC00003FFFFE00001FFFFF000007FFFF800003FFFFE00001FFFFF00000FFFFF800003FFFFE00001FFFFF000007FFFF800003FFFFE00000FFFFF000007FFFF";
defparam ram_block1a86.mem_init2 = "C00001FFFFE00000FFFFF800003FFFFE00001FFFFF000007FFFFC00001FFFFF000007FFFFC00003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800001FFFFF000007FFFFC00001FFFFF000003FFFFE00000FFFFF800003FFFFF000007FFFFC00001FFFFF800003FFFFE000007FFFFC00001FFFFF800003FFFFF000007FFFFE00000FFFFF800001FFFFF000003FFFFE000007FFFFE00000FFFFFC00001FFFFF800001FFFFF000003FFFFF000007FFFFE000007FFFFE00000FFFFFC00000FFFFFC00000FFFFF800001FFFFF800001FFFFF800001FFFFF800001FFFFF800001FFFFF";
defparam ram_block1a86.mem_init1 = "800001FFFFF800001FFFFF800001FFFFFC00000FFFFFC00000FFFFFC000007FFFFE000007FFFFF000003FFFFF000001FFFFF800000FFFFFC000007FFFFE000003FFFFF000001FFFFF800000FFFFFE000007FFFFF000001FFFFF800000FFFFFE000003FFFFF800001FFFFFC000007FFFFF000001FFFFFC000007FFFFF000001FFFFFC000003FFFFF800000FFFFFE000003FFFFFC000007FFFFF000000FFFFFE000003FFFFFC000007FFFFF800000FFFFFF000000FFFFFE000001FFFFFE000003FFFFFC000003FFFFFC000007FFFFF8000007FFFFF8000007FFFFF8000007FFFFF8000003FFFFFC000003FFFFFC000003FFFFFE000001FFFFFF000000FFFFFF000";
defparam ram_block1a86.mem_init0 = "0007FFFFF8000003FFFFFE000001FFFFFF0000007FFFFFC000003FFFFFE000000FFFFFF8000003FFFFFE000000FFFFFF8000003FFFFFF0000007FFFFFC000000FFFFFF8000003FFFFFF0000007FFFFFE0000007FFFFFC000000FFFFFFC000000FFFFFF8000001FFFFFF8000001FFFFFF8000000FFFFFFC000000FFFFFFC0000007FFFFFE0000007FFFFFF0000003FFFFFF8000000FFFFFFC0000007FFFFFF0000001FFFFFFC0000007FFFFFF0000001FFFFFFC0000003FFFFFF8000000FFFFFFF0000001FFFFFFE0000001FFFFFFE0000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000001FFFFFFE0000001FFFFFFF0000000FFFFFFF80000003FFFFFFC";

cyclonev_ram_block ram_block1a14(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "rom";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "clock0";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 8191;
defparam ram_block1a14.port_a_logical_ram_depth = 65536;
defparam ram_block1a14.port_a_logical_ram_width = 24;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init3 = "7FFFFFF80000003FFFFFFE0000001FFFFFFF0000000FFFFFFF00000007FFFFFF80000007FFFFFF80000007FFFFFF8000000FFFFFFF0000000FFFFFFF0000001FFFFFFE0000003FFFFFF80000007FFFFFF0000001FFFFFFC0000007FFFFFF0000001FFFFFFC0000007FFFFFE0000003FFFFFF8000001FFFFFFC000000FFFFFFC0000007FFFFFE0000007FFFFFE0000003FFFFFF0000003FFFFFF0000003FFFFFE0000007FFFFFE0000007FFFFFC000000FFFFFFC000001FFFFFF8000003FFFFFE0000007FFFFFC000001FFFFFF8000003FFFFFE000000FFFFFF8000003FFFFFE000000FFFFFF8000007FFFFFC000001FFFFFF000000FFFFFF8000003FFFFFC000";
defparam ram_block1a14.mem_init2 = "001FFFFFE000001FFFFFF000000FFFFFF8000007FFFFF8000007FFFFF8000003FFFFFC000003FFFFFC000003FFFFFC000003FFFFFC000007FFFFF8000007FFFFF800000FFFFFF000000FFFFFE000001FFFFFE000003FFFFFC000007FFFFF800000FFFFFE000001FFFFFC000007FFFFF800000FFFFFE000003FFFFF8000007FFFFF000001FFFFFC000007FFFFF000001FFFFFC000007FFFFF000003FFFFF800000FFFFFE000003FFFFF000001FFFFFC00000FFFFFE000003FFFFF000001FFFFF800000FFFFFC000007FFFFE000003FFFFF000001FFFFF800001FFFFFC00000FFFFFC000007FFFFE000007FFFFE000007FFFFF000003FFFFF000003FFFFF000003";
defparam ram_block1a14.mem_init1 = "FFFFF000003FFFFF000003FFFFF000003FFFFF000003FFFFF000003FFFFE000007FFFFE000007FFFFE00000FFFFFC00000FFFFFC00001FFFFF800001FFFFF000003FFFFF000007FFFFE00000FFFFFC00000FFFFF800001FFFFF000003FFFFE00000FFFFFC00001FFFFF800003FFFFF000007FFFFC00000FFFFF800003FFFFF000007FFFFC00001FFFFF800003FFFFE00000FFFFF800001FFFFF000007FFFFC00001FFFFF000003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800007FFFFC00001FFFFF000007FFFFC00001FFFFF00000FFFFF800003FFFFE00000FFFFF000007";
defparam ram_block1a14.mem_init0 = "FFFFC00001FFFFE00000FFFFF800003FFFFC00001FFFFF00000FFFFF800003FFFFE00001FFFFF00000FFFFF800003FFFFC00001FFFFF00000FFFFF800007FFFFC00001FFFFE00000FFFFF000007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFC00001FFFFE00000FFFFF000007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800007FFFFC00003FFFFE00001FFFFE00000FFFFF000007FFFF800007FFFFC00003FFFFC00001FFFFE00000";

cyclonev_ram_block ram_block1a38(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a38_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a38.clk0_core_clock_enable = "ena0";
defparam ram_block1a38.clk0_input_clock_enable = "ena0";
defparam ram_block1a38.clk0_output_clock_enable = "ena0";
defparam ram_block1a38.data_interleave_offset_in_bits = 1;
defparam ram_block1a38.data_interleave_width_in_bits = 1;
defparam ram_block1a38.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a38.init_file_layout = "port_a";
defparam ram_block1a38.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a38.operation_mode = "rom";
defparam ram_block1a38.port_a_address_clear = "none";
defparam ram_block1a38.port_a_address_width = 13;
defparam ram_block1a38.port_a_data_out_clear = "none";
defparam ram_block1a38.port_a_data_out_clock = "clock0";
defparam ram_block1a38.port_a_data_width = 1;
defparam ram_block1a38.port_a_first_address = 8192;
defparam ram_block1a38.port_a_first_bit_number = 14;
defparam ram_block1a38.port_a_last_address = 16383;
defparam ram_block1a38.port_a_logical_ram_depth = 65536;
defparam ram_block1a38.port_a_logical_ram_width = 24;
defparam ram_block1a38.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a38.ram_block_type = "auto";
defparam ram_block1a38.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000";
defparam ram_block1a38.mem_init2 = "0000FFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFFFFFFFFFC000000000000000000003FFFFFFFFFFFFFFFFFFFE00000000000000000007FFFFFFFFFFFFFFFFFFC000000000000000000FFFFFFFFFFFFFFFFFF800000000000000000FFFFFFFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFF00000000000000003FFFFFFFFFFFFFFFC0000000000000007FFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFF000000000000001FFFFFFFFFFFFFF800000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFF80000000000001FFFFFFFFFFFFF";
defparam ram_block1a38.mem_init1 = "80000000000003FFFFFFFFFFFFC0000000000003FFFFFFFFFFFF8000000000001FFFFFFFFFFFF8000000000001FFFFFFFFFFFF000000000000FFFFFFFFFFFF000000000001FFFFFFFFFFFE000000000007FFFFFFFFFFE000000000007FFFFFFFFFFC00000000001FFFFFFFFFFF00000000000FFFFFFFFFFF00000000000FFFFFFFFFFE00000000003FFFFFFFFFF00000000001FFFFFFFFFF80000000003FFFFFFFFFE00000000007FFFFFFFFF80000000003FFFFFFFFFC0000000003FFFFFFFFFC0000000007FFFFFFFFF0000000001FFFFFFFFFC0000000007FFFFFFFFE0000000007FFFFFFFFE000000000FFFFFFFFFC000000001FFFFFFFFF0000000007FF";
defparam ram_block1a38.mem_init0 = "FFFFFFC000000003FFFFFFFFC000000003FFFFFFFFC000000003FFFFFFFF8000000007FFFFFFFF000000001FFFFFFFFC000000007FFFFFFFE000000003FFFFFFFF000000003FFFFFFFF000000003FFFFFFFE000000007FFFFFFFC00000001FFFFFFFF000000007FFFFFFFC00000001FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF800000007FFFFFFF00000000FFFFFFFF00000001FFFFFFFE00000003FFFFFFF80000000FFFFFFFE00000003FFFFFFF80000001FFFFFFFC0000000FFFFFFFE00000007FFFFFFE00000007FFFFFFE00000007FFFFFFE0000000FFFFFFFC0000000FFFFFFF80000003FFFFFFF00000007FFFFFFC0000001FFFFFFF0000000";

cyclonev_ram_block ram_block1a111(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a111_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a111.clk0_core_clock_enable = "ena0";
defparam ram_block1a111.clk0_input_clock_enable = "ena0";
defparam ram_block1a111.clk0_output_clock_enable = "ena0";
defparam ram_block1a111.data_interleave_offset_in_bits = 1;
defparam ram_block1a111.data_interleave_width_in_bits = 1;
defparam ram_block1a111.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a111.init_file_layout = "port_a";
defparam ram_block1a111.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a111.operation_mode = "rom";
defparam ram_block1a111.port_a_address_clear = "none";
defparam ram_block1a111.port_a_address_width = 13;
defparam ram_block1a111.port_a_data_out_clear = "none";
defparam ram_block1a111.port_a_data_out_clock = "clock0";
defparam ram_block1a111.port_a_data_width = 1;
defparam ram_block1a111.port_a_first_address = 32768;
defparam ram_block1a111.port_a_first_bit_number = 15;
defparam ram_block1a111.port_a_last_address = 40959;
defparam ram_block1a111.port_a_logical_ram_depth = 65536;
defparam ram_block1a111.port_a_logical_ram_width = 24;
defparam ram_block1a111.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a111.ram_block_type = "auto";
defparam ram_block1a111.mem_init3 = "7FFFFFFFFFFFFFC00000000000001FFFFFFFFFFFFFF000000000000007FFFFFFFFFFFFF800000000000007FFFFFFFFFFFFF00000000000000FFFFFFFFFFFFFE00000000000003FFFFFFFFFFFFF80000000000001FFFFFFFFFFFFF80000000000001FFFFFFFFFFFFF80000000000003FFFFFFFFFFFFE0000000000000FFFFFFFFFFFFF80000000000007FFFFFFFFFFFFC0000000000003FFFFFFFFFFFFC0000000000007FFFFFFFFFFFF8000000000000FFFFFFFFFFFFE0000000000003FFFFFFFFFFFF8000000000001FFFFFFFFFFFFC000000000000FFFFFFFFFFFFC000000000000FFFFFFFFFFFF8000000000001FFFFFFFFFFFF0000000000003FFFFFFFFF";
defparam ram_block1a111.mem_init2 = "FFE000000000001FFFFFFFFFFFF0000000000007FFFFFFFFFFF8000000000003FFFFFFFFFFFC000000000003FFFFFFFFFFFC000000000007FFFFFFFFFFF800000000000FFFFFFFFFFFF000000000001FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000001FFFFFFFFFFF800000000000FFFFFFFFFFFC000000000007FFFFFFFFFFE000000000007FFFFFFFFFFE000000000007FFFFFFFFFFC00000000000FFFFFFFFFFFC00000000001FFFFFFFFFFF000000000003FFFFFFFFFFE00000000000FFFFFFFFFFF800000000003FFFFFFFFFFE00000000001FFFFFFFFFFF000000000007FFFFFFFFFF800000000007FFFFFFFFFFC00000000003FFFFFFFFFFC";
defparam ram_block1a111.mem_init1 = "00000000003FFFFFFFFFFC00000000003FFFFFFFFFFC00000000003FFFFFFFFFF800000000007FFFFFFFFFF00000000000FFFFFFFFFFE00000000001FFFFFFFFFFC00000000007FFFFFFFFFF00000000000FFFFFFFFFFE00000000003FFFFFFFFFF00000000001FFFFFFFFFFC00000000007FFFFFFFFFF00000000003FFFFFFFFFF80000000001FFFFFFFFFFC0000000000FFFFFFFFFFE00000000007FFFFFFFFFE00000000003FFFFFFFFFF00000000003FFFFFFFFFF00000000003FFFFFFFFFF00000000003FFFFFFFFFF00000000003FFFFFFFFFF00000000007FFFFFFFFFE00000000007FFFFFFFFFE0000000000FFFFFFFFFFC0000000000FFFFFFFFFF8";
defparam ram_block1a111.mem_init0 = "0000000001FFFFFFFFFF00000000003FFFFFFFFFE0000000000FFFFFFFFFFC0000000001FFFFFFFFFF00000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000007FFFFFFFFFC0000000001FFFFFFFFFE";

cyclonev_ram_block ram_block1a135(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a135_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a135.clk0_core_clock_enable = "ena0";
defparam ram_block1a135.clk0_input_clock_enable = "ena0";
defparam ram_block1a135.clk0_output_clock_enable = "ena0";
defparam ram_block1a135.data_interleave_offset_in_bits = 1;
defparam ram_block1a135.data_interleave_width_in_bits = 1;
defparam ram_block1a135.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a135.init_file_layout = "port_a";
defparam ram_block1a135.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a135.operation_mode = "rom";
defparam ram_block1a135.port_a_address_clear = "none";
defparam ram_block1a135.port_a_address_width = 13;
defparam ram_block1a135.port_a_data_out_clear = "none";
defparam ram_block1a135.port_a_data_out_clock = "clock0";
defparam ram_block1a135.port_a_data_width = 1;
defparam ram_block1a135.port_a_first_address = 40960;
defparam ram_block1a135.port_a_first_bit_number = 15;
defparam ram_block1a135.port_a_last_address = 49151;
defparam ram_block1a135.port_a_logical_ram_depth = 65536;
defparam ram_block1a135.port_a_logical_ram_width = 24;
defparam ram_block1a135.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a135.ram_block_type = "auto";
defparam ram_block1a135.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000";
defparam ram_block1a135.mem_init2 = "0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000001FFFFFFFFFFFFF";
defparam ram_block1a135.mem_init1 = "FFFFFFFFFFFFFC00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000007FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFFFFFFFFFE000000000000000000003FFFFFFFFFFFFFFFFFFFF800000000000000000003FFFFFFFFFFFFFFFFFFFC00000000000000000007FFFFFFFFFFFFFFFFFFE00000000000000000007FFFFFFFFFFFFFFFFFF8000000000000000000FFFFFFFFFFFFFFFFFFE0000000000000000007FF";
defparam ram_block1a135.mem_init0 = "FFFFFFFFFFFFFFFC000000000000000003FFFFFFFFFFFFFFFFFC000000000000000007FFFFFFFFFFFFFFFFE000000000000000007FFFFFFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFFC00000000000000007FFFFFFFFFFFFFFFE00000000000000007FFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFFFFFF00000000000000007FFFFFFFFFFFFFFF0000000000000001FFFFFFFFFFFFFFFC000000000000000FFFFFFFFFFFFFFFC000000000000001FFFFFFFFFFFFFFF0000000000000007FFFFFFFFFFFFFF8000000000000007FFFFFFFFFFFFFF000000000000000FFFFFFFFFFFFFFC000000000000007FFFFFFFFFFFFFE00000000000000";

cyclonev_ram_block ram_block1a159(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a159_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a159.clk0_core_clock_enable = "ena0";
defparam ram_block1a159.clk0_input_clock_enable = "ena0";
defparam ram_block1a159.clk0_output_clock_enable = "ena0";
defparam ram_block1a159.data_interleave_offset_in_bits = 1;
defparam ram_block1a159.data_interleave_width_in_bits = 1;
defparam ram_block1a159.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a159.init_file_layout = "port_a";
defparam ram_block1a159.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a159.operation_mode = "rom";
defparam ram_block1a159.port_a_address_clear = "none";
defparam ram_block1a159.port_a_address_width = 13;
defparam ram_block1a159.port_a_data_out_clear = "none";
defparam ram_block1a159.port_a_data_out_clock = "clock0";
defparam ram_block1a159.port_a_data_width = 1;
defparam ram_block1a159.port_a_first_address = 49152;
defparam ram_block1a159.port_a_first_bit_number = 15;
defparam ram_block1a159.port_a_last_address = 57343;
defparam ram_block1a159.port_a_logical_ram_depth = 65536;
defparam ram_block1a159.port_a_logical_ram_width = 24;
defparam ram_block1a159.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a159.ram_block_type = "auto";
defparam ram_block1a159.mem_init3 = "00000000000000FFFFFFFFFFFFFFC000000000000007FFFFFFFFFFFFFE000000000000001FFFFFFFFFFFFFFC000000000000003FFFFFFFFFFFFFFC000000000000001FFFFFFFFFFFFFFF0000000000000007FFFFFFFFFFFFFFE0000000000000007FFFFFFFFFFFFFFF0000000000000001FFFFFFFFFFFFFFFC0000000000000001FFFFFFFFFFFFFFFE0000000000000000FFFFFFFFFFFFFFFFC0000000000000000FFFFFFFFFFFFFFFFC00000000000000007FFFFFFFFFFFFFFFF800000000000000007FFFFFFFFFFFFFFFFC00000000000000000FFFFFFFFFFFFFFFFFC000000000000000007FFFFFFFFFFFFFFFFF8000000000000000007FFFFFFFFFFFFFFF";
defparam ram_block1a159.mem_init2 = "FFC000000000000000000FFFFFFFFFFFFFFFFFFE0000000000000000003FFFFFFFFFFFFFFFFFFC0000000000000000000FFFFFFFFFFFFFFFFFFFC00000000000000000007FFFFFFFFFFFFFFFFFFF800000000000000000003FFFFFFFFFFFFFFFFFFFF800000000000000000000FFFFFFFFFFFFFFFFFFFFF8000000000000000000001FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000007FFFFFFFFFFFFF";
defparam ram_block1a159.mem_init1 = "FFFFFFFFFFFFF0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000";
defparam ram_block1a159.mem_init0 = "000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a183(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a183_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a183.clk0_core_clock_enable = "ena0";
defparam ram_block1a183.clk0_input_clock_enable = "ena0";
defparam ram_block1a183.clk0_output_clock_enable = "ena0";
defparam ram_block1a183.data_interleave_offset_in_bits = 1;
defparam ram_block1a183.data_interleave_width_in_bits = 1;
defparam ram_block1a183.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a183.init_file_layout = "port_a";
defparam ram_block1a183.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a183.operation_mode = "rom";
defparam ram_block1a183.port_a_address_clear = "none";
defparam ram_block1a183.port_a_address_width = 13;
defparam ram_block1a183.port_a_data_out_clear = "none";
defparam ram_block1a183.port_a_data_out_clock = "clock0";
defparam ram_block1a183.port_a_data_width = 1;
defparam ram_block1a183.port_a_first_address = 57344;
defparam ram_block1a183.port_a_first_bit_number = 15;
defparam ram_block1a183.port_a_last_address = 65535;
defparam ram_block1a183.port_a_logical_ram_depth = 65536;
defparam ram_block1a183.port_a_logical_ram_width = 24;
defparam ram_block1a183.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a183.ram_block_type = "auto";
defparam ram_block1a183.mem_init3 = "FFFFFFFFFF00000000007FFFFFFFFFC0000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000001FFFFFFFFFF00000000007FFFFFFFFFE0000000000FFFFFFFFFF80000000001FFFFFFFFFF0000000000";
defparam ram_block1a183.mem_init2 = "3FFFFFFFFFE00000000007FFFFFFFFFE0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000001FFFFFFFFFF80000000001FFFFFFFFFF80000000001FFFFFFFFFF80000000001FFFFFFFFFF80000000001FFFFFFFFFF80000000000FFFFFFFFFFC0000000000FFFFFFFFFFE00000000007FFFFFFFFFF00000000003FFFFFFFFFF80000000001FFFFFFFFFFC00000000007FFFFFFFFFF00000000001FFFFFFFFFF80000000000FFFFFFFFFFE00000000001FFFFFFFFFFC00000000007FFFFFFFFFF00000000000FFFFFFFFFFE00000000001FFFFFFFFFFC00000000003FFFFFFFFFF800000000007FFFFFFFFFF800000000007FFFFFFFFFF80000000000";
defparam ram_block1a183.mem_init1 = "7FFFFFFFFFF800000000007FFFFFFFFFFC00000000003FFFFFFFFFFC00000000001FFFFFFFFFFF00000000000FFFFFFFFFFF800000000003FFFFFFFFFFE00000000000FFFFFFFFFFF800000000001FFFFFFFFFFF000000000007FFFFFFFFFFE000000000007FFFFFFFFFFC00000000000FFFFFFFFFFFC00000000000FFFFFFFFFFFC000000000007FFFFFFFFFFE000000000003FFFFFFFFFFF000000000001FFFFFFFFFFFC000000000007FFFFFFFFFFF000000000001FFFFFFFFFFFE000000000003FFFFFFFFFFFC000000000007FFFFFFFFFFF8000000000007FFFFFFFFFFF8000000000003FFFFFFFFFFFC000000000001FFFFFFFFFFFF000000000000FFF";
defparam ram_block1a183.mem_init0 = "FFFFFFFFF8000000000001FFFFFFFFFFFF0000000000003FFFFFFFFFFFE0000000000007FFFFFFFFFFFE0000000000007FFFFFFFFFFFF0000000000003FFFFFFFFFFFF8000000000000FFFFFFFFFFFFE0000000000003FFFFFFFFFFFFC0000000000007FFFFFFFFFFFF80000000000007FFFFFFFFFFFFC0000000000003FFFFFFFFFFFFE0000000000000FFFFFFFFFFFFF80000000000003FFFFFFFFFFFFF00000000000003FFFFFFFFFFFFF00000000000003FFFFFFFFFFFFF80000000000000FFFFFFFFFFFFFE00000000000001FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFC00000000000001FFFFFFFFFFFFFF000000000000007FFFFFFFFFFFFFC";

cyclonev_ram_block ram_block1a63(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a63_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a63.clk0_core_clock_enable = "ena0";
defparam ram_block1a63.clk0_input_clock_enable = "ena0";
defparam ram_block1a63.clk0_output_clock_enable = "ena0";
defparam ram_block1a63.data_interleave_offset_in_bits = 1;
defparam ram_block1a63.data_interleave_width_in_bits = 1;
defparam ram_block1a63.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a63.init_file_layout = "port_a";
defparam ram_block1a63.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a63.operation_mode = "rom";
defparam ram_block1a63.port_a_address_clear = "none";
defparam ram_block1a63.port_a_address_width = 13;
defparam ram_block1a63.port_a_data_out_clear = "none";
defparam ram_block1a63.port_a_data_out_clock = "clock0";
defparam ram_block1a63.port_a_data_width = 1;
defparam ram_block1a63.port_a_first_address = 16384;
defparam ram_block1a63.port_a_first_bit_number = 15;
defparam ram_block1a63.port_a_last_address = 24575;
defparam ram_block1a63.port_a_logical_ram_depth = 65536;
defparam ram_block1a63.port_a_logical_ram_width = 24;
defparam ram_block1a63.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a63.ram_block_type = "auto";
defparam ram_block1a63.mem_init3 = "FFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFF800000000000001FFFFFFFFFFFFFFE000000000000003FFFFFFFFFFFFFFC000000000000003FFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFF8000000000000001FFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFE0000000000000003FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFFF00000000000000003FFFFFFFFFFFFFFFF00000000000000003FFFFFFFFFFFFFFFF800000000000000007FFFFFFFFFFFFFFFF800000000000000003FFFFFFFFFFFFFFFFF000000000000000003FFFFFFFFFFFFFFFFF8000000000000000007FFFFFFFFFFFFFFFFF8000000000000000";
defparam ram_block1a63.mem_init2 = "003FFFFFFFFFFFFFFFFFF0000000000000000001FFFFFFFFFFFFFFFFFFC0000000000000000003FFFFFFFFFFFFFFFFFFF00000000000000000003FFFFFFFFFFFFFFFFFFF800000000000000000007FFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFF0000000000000000000007FFFFFFFFFFFFFFFFFFFFE0000000000000000000001FFFFFFFFFFFFFFFFFFFFFF00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF80000000000000";
defparam ram_block1a63.mem_init1 = "0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000001FFFF";
defparam ram_block1a63.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a87(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a87_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a87.clk0_core_clock_enable = "ena0";
defparam ram_block1a87.clk0_input_clock_enable = "ena0";
defparam ram_block1a87.clk0_output_clock_enable = "ena0";
defparam ram_block1a87.data_interleave_offset_in_bits = 1;
defparam ram_block1a87.data_interleave_width_in_bits = 1;
defparam ram_block1a87.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a87.init_file_layout = "port_a";
defparam ram_block1a87.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a87.operation_mode = "rom";
defparam ram_block1a87.port_a_address_clear = "none";
defparam ram_block1a87.port_a_address_width = 13;
defparam ram_block1a87.port_a_data_out_clear = "none";
defparam ram_block1a87.port_a_data_out_clock = "clock0";
defparam ram_block1a87.port_a_data_width = 1;
defparam ram_block1a87.port_a_first_address = 24576;
defparam ram_block1a87.port_a_first_bit_number = 15;
defparam ram_block1a87.port_a_last_address = 32767;
defparam ram_block1a87.port_a_logical_ram_depth = 65536;
defparam ram_block1a87.port_a_logical_ram_width = 24;
defparam ram_block1a87.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a87.ram_block_type = "auto";
defparam ram_block1a87.mem_init3 = "0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFE0000000000FFFFFFFFFF80000000001FFFFFFFFFF00000000007FFFFFFFFFE0000000000FFFFFFFFFF";
defparam ram_block1a87.mem_init2 = "C0000000001FFFFFFFFFF80000000001FFFFFFFFFF00000000003FFFFFFFFFF00000000003FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFF00000000003FFFFFFFFFF00000000001FFFFFFFFFF80000000000FFFFFFFFFFC00000000007FFFFFFFFFE00000000003FFFFFFFFFF80000000000FFFFFFFFFFE00000000007FFFFFFFFFF00000000001FFFFFFFFFFE00000000003FFFFFFFFFF80000000000FFFFFFFFFFF00000000001FFFFFFFFFFE00000000003FFFFFFFFFFC00000000007FFFFFFFFFF800000000007FFFFFFFFFF800000000007FFFFFFFFFF";
defparam ram_block1a87.mem_init1 = "800000000007FFFFFFFFFF800000000003FFFFFFFFFFC00000000003FFFFFFFFFFE00000000000FFFFFFFFFFF000000000007FFFFFFFFFFC00000000001FFFFFFFFFFF000000000007FFFFFFFFFFE00000000000FFFFFFFFFFF800000000001FFFFFFFFFFF800000000003FFFFFFFFFFF000000000003FFFFFFFFFFF000000000003FFFFFFFFFFF800000000001FFFFFFFFFFFC00000000000FFFFFFFFFFFE000000000003FFFFFFFFFFF800000000000FFFFFFFFFFFE000000000001FFFFFFFFFFFC000000000003FFFFFFFFFFF8000000000007FFFFFFFFFFF8000000000007FFFFFFFFFFFC000000000003FFFFFFFFFFFE000000000000FFFFFFFFFFFF000";
defparam ram_block1a87.mem_init0 = "0000000007FFFFFFFFFFFE000000000000FFFFFFFFFFFFC000000000001FFFFFFFFFFFF8000000000001FFFFFFFFFFFF8000000000000FFFFFFFFFFFFC0000000000007FFFFFFFFFFFF0000000000001FFFFFFFFFFFFC0000000000003FFFFFFFFFFFF80000000000007FFFFFFFFFFFF80000000000003FFFFFFFFFFFFC0000000000001FFFFFFFFFFFFF00000000000007FFFFFFFFFFFFC0000000000000FFFFFFFFFFFFFC0000000000000FFFFFFFFFFFFFC00000000000007FFFFFFFFFFFFF00000000000001FFFFFFFFFFFFFE00000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFE00000000000000FFFFFFFFFFFFFF800000000000003";

cyclonev_ram_block ram_block1a15(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "rom";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "clock0";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 8191;
defparam ram_block1a15.port_a_logical_ram_depth = 65536;
defparam ram_block1a15.port_a_logical_ram_width = 24;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init3 = "800000000000003FFFFFFFFFFFFFE00000000000000FFFFFFFFFFFFFF800000000000007FFFFFFFFFFFFF80000000000000FFFFFFFFFFFFFF00000000000001FFFFFFFFFFFFFC00000000000007FFFFFFFFFFFFE00000000000007FFFFFFFFFFFFE00000000000007FFFFFFFFFFFFC0000000000001FFFFFFFFFFFFF00000000000007FFFFFFFFFFFF80000000000003FFFFFFFFFFFFC0000000000003FFFFFFFFFFFF80000000000007FFFFFFFFFFFF0000000000001FFFFFFFFFFFFC0000000000007FFFFFFFFFFFE0000000000003FFFFFFFFFFFF0000000000003FFFFFFFFFFFF0000000000007FFFFFFFFFFFE000000000000FFFFFFFFFFFFC000000000";
defparam ram_block1a15.mem_init2 = "001FFFFFFFFFFFE000000000000FFFFFFFFFFFF8000000000007FFFFFFFFFFFC000000000003FFFFFFFFFFFC000000000003FFFFFFFFFFF8000000000007FFFFFFFFFFF000000000000FFFFFFFFFFFE000000000003FFFFFFFFFFF800000000000FFFFFFFFFFFE000000000007FFFFFFFFFFF000000000003FFFFFFFFFFF800000000001FFFFFFFFFFF800000000001FFFFFFFFFFF800000000003FFFFFFFFFFF000000000003FFFFFFFFFFE00000000000FFFFFFFFFFFC00000000001FFFFFFFFFFF000000000007FFFFFFFFFFC00000000001FFFFFFFFFFE00000000000FFFFFFFFFFF800000000007FFFFFFFFFF800000000003FFFFFFFFFFC00000000003";
defparam ram_block1a15.mem_init1 = "FFFFFFFFFFC00000000003FFFFFFFFFFC00000000003FFFFFFFFFFC00000000007FFFFFFFFFF80000000000FFFFFFFFFFF00000000001FFFFFFFFFFE00000000003FFFFFFFFFF80000000000FFFFFFFFFFF00000000001FFFFFFFFFFC0000000000FFFFFFFFFFE00000000003FFFFFFFFFF80000000000FFFFFFFFFFC00000000007FFFFFFFFFE00000000003FFFFFFFFFF00000000001FFFFFFFFFF80000000001FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFF80000000001FFFFFFFFFF80000000001FFFFFFFFFF00000000003FFFFFFFFFF00000000007";
defparam ram_block1a15.mem_init0 = "FFFFFFFFFE0000000000FFFFFFFFFFC0000000001FFFFFFFFFF00000000003FFFFFFFFFE0000000000FFFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFE0000000000";

cyclonev_ram_block ram_block1a39(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a39_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a39.clk0_core_clock_enable = "ena0";
defparam ram_block1a39.clk0_input_clock_enable = "ena0";
defparam ram_block1a39.clk0_output_clock_enable = "ena0";
defparam ram_block1a39.data_interleave_offset_in_bits = 1;
defparam ram_block1a39.data_interleave_width_in_bits = 1;
defparam ram_block1a39.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a39.init_file_layout = "port_a";
defparam ram_block1a39.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a39.operation_mode = "rom";
defparam ram_block1a39.port_a_address_clear = "none";
defparam ram_block1a39.port_a_address_width = 13;
defparam ram_block1a39.port_a_data_out_clear = "none";
defparam ram_block1a39.port_a_data_out_clock = "clock0";
defparam ram_block1a39.port_a_data_width = 1;
defparam ram_block1a39.port_a_first_address = 8192;
defparam ram_block1a39.port_a_first_bit_number = 15;
defparam ram_block1a39.port_a_last_address = 16383;
defparam ram_block1a39.port_a_logical_ram_depth = 65536;
defparam ram_block1a39.port_a_logical_ram_width = 24;
defparam ram_block1a39.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a39.ram_block_type = "auto";
defparam ram_block1a39.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a39.mem_init2 = "FFFF00000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000";
defparam ram_block1a39.mem_init1 = "00000000000003FFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000007FFFFFFFFFFFFFFFFFFFFFF80000000000000000000001FFFFFFFFFFFFFFFFFFFFFF0000000000000000000000FFFFFFFFFFFFFFFFFFFFFC000000000000000000001FFFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000003FFFFFFFFFFFFFFFFFFF80000000000000000001FFFFFFFFFFFFFFFFFFF80000000000000000007FFFFFFFFFFFFFFFFFF0000000000000000001FFFFFFFFFFFFFFFFFF800";
defparam ram_block1a39.mem_init0 = "0000000000000003FFFFFFFFFFFFFFFFFC000000000000000003FFFFFFFFFFFFFFFFF800000000000000001FFFFFFFFFFFFFFFFF800000000000000003FFFFFFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFF80000000000000001FFFFFFFFFFFFFFFF80000000000000001FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFE0000000000000003FFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFF8000000000000007FFFFFFFFFFFFFF800000000000000FFFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFF800000000000001FFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a112(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a112_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a112.clk0_core_clock_enable = "ena0";
defparam ram_block1a112.clk0_input_clock_enable = "ena0";
defparam ram_block1a112.clk0_output_clock_enable = "ena0";
defparam ram_block1a112.data_interleave_offset_in_bits = 1;
defparam ram_block1a112.data_interleave_width_in_bits = 1;
defparam ram_block1a112.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a112.init_file_layout = "port_a";
defparam ram_block1a112.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a112.operation_mode = "rom";
defparam ram_block1a112.port_a_address_clear = "none";
defparam ram_block1a112.port_a_address_width = 13;
defparam ram_block1a112.port_a_data_out_clear = "none";
defparam ram_block1a112.port_a_data_out_clock = "clock0";
defparam ram_block1a112.port_a_data_width = 1;
defparam ram_block1a112.port_a_first_address = 32768;
defparam ram_block1a112.port_a_first_bit_number = 16;
defparam ram_block1a112.port_a_last_address = 40959;
defparam ram_block1a112.port_a_logical_ram_depth = 65536;
defparam ram_block1a112.port_a_logical_ram_width = 24;
defparam ram_block1a112.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a112.ram_block_type = "auto";
defparam ram_block1a112.mem_init3 = "FFFFFFFFFFFFFFC0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000";
defparam ram_block1a112.mem_init2 = "001FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000003FFFFFFFFFFFFFFFFFFFFFFE00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000003FFFFFFFFFFFFFFFFFFFFFF00000000000000000000001FFFFFFFFFFFFFFFFFFFFFF80000000000000000000001FFFFFFFFFFFFFFFFFFFFFF00000000000000000000007FFFFFFFFFFFFFFFFFFFFFC0000000000000000000003";
defparam ram_block1a112.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC0000000000000000000003FFFFFFFFFFFFFFFFFFFFF8000000000000000000000FFFFFFFFFFFFFFFFFFFFFE0000000000000000000003FFFFFFFFFFFFFFFFFFFFF0000000000000000000001FFFFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFFFFFFFFFF0000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFC000000000000000000007";
defparam ram_block1a112.mem_init0 = "FFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000003FFFFFFFFFFFFFFFFFFFE";

cyclonev_ram_block ram_block1a136(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a136_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a136.clk0_core_clock_enable = "ena0";
defparam ram_block1a136.clk0_input_clock_enable = "ena0";
defparam ram_block1a136.clk0_output_clock_enable = "ena0";
defparam ram_block1a136.data_interleave_offset_in_bits = 1;
defparam ram_block1a136.data_interleave_width_in_bits = 1;
defparam ram_block1a136.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a136.init_file_layout = "port_a";
defparam ram_block1a136.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a136.operation_mode = "rom";
defparam ram_block1a136.port_a_address_clear = "none";
defparam ram_block1a136.port_a_address_width = 13;
defparam ram_block1a136.port_a_data_out_clear = "none";
defparam ram_block1a136.port_a_data_out_clock = "clock0";
defparam ram_block1a136.port_a_data_width = 1;
defparam ram_block1a136.port_a_first_address = 40960;
defparam ram_block1a136.port_a_first_bit_number = 16;
defparam ram_block1a136.port_a_last_address = 49151;
defparam ram_block1a136.port_a_logical_ram_depth = 65536;
defparam ram_block1a136.port_a_logical_ram_width = 24;
defparam ram_block1a136.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a136.ram_block_type = "auto";
defparam ram_block1a136.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000";
defparam ram_block1a136.mem_init2 = "000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a136.mem_init1 = "FFFFFFFFFFFFFC000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a136.mem_init0 = "FFFFFFFFFFFFFFFC000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000001FFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a160(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a160_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a160.clk0_core_clock_enable = "ena0";
defparam ram_block1a160.clk0_input_clock_enable = "ena0";
defparam ram_block1a160.clk0_output_clock_enable = "ena0";
defparam ram_block1a160.data_interleave_offset_in_bits = 1;
defparam ram_block1a160.data_interleave_width_in_bits = 1;
defparam ram_block1a160.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a160.init_file_layout = "port_a";
defparam ram_block1a160.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a160.operation_mode = "rom";
defparam ram_block1a160.port_a_address_clear = "none";
defparam ram_block1a160.port_a_address_width = 13;
defparam ram_block1a160.port_a_data_out_clear = "none";
defparam ram_block1a160.port_a_data_out_clock = "clock0";
defparam ram_block1a160.port_a_data_width = 1;
defparam ram_block1a160.port_a_first_address = 49152;
defparam ram_block1a160.port_a_first_bit_number = 16;
defparam ram_block1a160.port_a_last_address = 57343;
defparam ram_block1a160.port_a_logical_ram_depth = 65536;
defparam ram_block1a160.port_a_logical_ram_width = 24;
defparam ram_block1a160.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a160.ram_block_type = "auto";
defparam ram_block1a160.mem_init3 = "FFFFFFFFFFFFFF000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000007FFFFFFFFFFFFFFF";
defparam ram_block1a160.mem_init2 = "FFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000007FFFFFFFFFFFFF";
defparam ram_block1a160.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000";
defparam ram_block1a160.mem_init0 = "000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a184(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a184_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a184.clk0_core_clock_enable = "ena0";
defparam ram_block1a184.clk0_input_clock_enable = "ena0";
defparam ram_block1a184.clk0_output_clock_enable = "ena0";
defparam ram_block1a184.data_interleave_offset_in_bits = 1;
defparam ram_block1a184.data_interleave_width_in_bits = 1;
defparam ram_block1a184.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a184.init_file_layout = "port_a";
defparam ram_block1a184.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a184.operation_mode = "rom";
defparam ram_block1a184.port_a_address_clear = "none";
defparam ram_block1a184.port_a_address_width = 13;
defparam ram_block1a184.port_a_data_out_clear = "none";
defparam ram_block1a184.port_a_data_out_clock = "clock0";
defparam ram_block1a184.port_a_data_width = 1;
defparam ram_block1a184.port_a_first_address = 57344;
defparam ram_block1a184.port_a_first_bit_number = 16;
defparam ram_block1a184.port_a_last_address = 65535;
defparam ram_block1a184.port_a_logical_ram_depth = 65536;
defparam ram_block1a184.port_a_logical_ram_width = 24;
defparam ram_block1a184.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a184.ram_block_type = "auto";
defparam ram_block1a184.mem_init3 = "FFFFFFFFFFFFFFFFFFFF800000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a184.mem_init2 = "C000000000000000000007FFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000000FFFFFFFFFFFFFFFFFFFFF0000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000001FFFFFFFFFFFFFFFFFFFFF8000000000000000000001FFFFFFFFFFFFFFFFFFFFF0000000000000000000001FFFFFFFFFFFFFFFFFFFFF8000000000000000000000FFFFFFFFFFFFFFFFFFFFFE0000000000000000000003FFFFFFFFFFFFFFFFFFFFF80000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a184.mem_init1 = "80000000000000000000007FFFFFFFFFFFFFFFFFFFFFC0000000000000000000001FFFFFFFFFFFFFFFFFFFFFF00000000000000000000003FFFFFFFFFFFFFFFFFFFFFF00000000000000000000001FFFFFFFFFFFFFFFFFFFFFF800000000000000000000007FFFFFFFFFFFFFFFFFFFFFF00000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000003FFFFFFFFFFFFFFFFFFFFFFE000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFE000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFF000";
defparam ram_block1a184.mem_init0 = "0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000007FFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a64(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a64_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a64.clk0_core_clock_enable = "ena0";
defparam ram_block1a64.clk0_input_clock_enable = "ena0";
defparam ram_block1a64.clk0_output_clock_enable = "ena0";
defparam ram_block1a64.data_interleave_offset_in_bits = 1;
defparam ram_block1a64.data_interleave_width_in_bits = 1;
defparam ram_block1a64.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a64.init_file_layout = "port_a";
defparam ram_block1a64.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a64.operation_mode = "rom";
defparam ram_block1a64.port_a_address_clear = "none";
defparam ram_block1a64.port_a_address_width = 13;
defparam ram_block1a64.port_a_data_out_clear = "none";
defparam ram_block1a64.port_a_data_out_clock = "clock0";
defparam ram_block1a64.port_a_data_width = 1;
defparam ram_block1a64.port_a_first_address = 16384;
defparam ram_block1a64.port_a_first_bit_number = 16;
defparam ram_block1a64.port_a_last_address = 24575;
defparam ram_block1a64.port_a_logical_ram_depth = 65536;
defparam ram_block1a64.port_a_logical_ram_width = 24;
defparam ram_block1a64.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a64.ram_block_type = "auto";
defparam ram_block1a64.mem_init3 = "00000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000";
defparam ram_block1a64.mem_init2 = "000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000";
defparam ram_block1a64.mem_init1 = "00000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a64.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a88(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a88_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a88.clk0_core_clock_enable = "ena0";
defparam ram_block1a88.clk0_input_clock_enable = "ena0";
defparam ram_block1a88.clk0_output_clock_enable = "ena0";
defparam ram_block1a88.data_interleave_offset_in_bits = 1;
defparam ram_block1a88.data_interleave_width_in_bits = 1;
defparam ram_block1a88.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a88.init_file_layout = "port_a";
defparam ram_block1a88.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a88.operation_mode = "rom";
defparam ram_block1a88.port_a_address_clear = "none";
defparam ram_block1a88.port_a_address_width = 13;
defparam ram_block1a88.port_a_data_out_clear = "none";
defparam ram_block1a88.port_a_data_out_clock = "clock0";
defparam ram_block1a88.port_a_data_width = 1;
defparam ram_block1a88.port_a_first_address = 24576;
defparam ram_block1a88.port_a_first_bit_number = 16;
defparam ram_block1a88.port_a_last_address = 32767;
defparam ram_block1a88.port_a_logical_ram_depth = 65536;
defparam ram_block1a88.port_a_logical_ram_width = 24;
defparam ram_block1a88.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a88.ram_block_type = "auto";
defparam ram_block1a88.mem_init3 = "000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000000FFFFFFFFFFFFFFFFFFFFE00000000000000000000";
defparam ram_block1a88.mem_init2 = "3FFFFFFFFFFFFFFFFFFFF800000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF8000000000000000000003FFFFFFFFFFFFFFFFFFFFE0000000000000000000007FFFFFFFFFFFFFFFFFFFFE000000000000000000000FFFFFFFFFFFFFFFFFFFFFE0000000000000000000007FFFFFFFFFFFFFFFFFFFFF0000000000000000000001FFFFFFFFFFFFFFFFFFFFFC0000000000000000000007FFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a88.mem_init1 = "7FFFFFFFFFFFFFFFFFFFFF80000000000000000000003FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFE00000000000000000000007FFFFFFFFFFFFFFFFFFFFFF80000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF800000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000FFF";
defparam ram_block1a88.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000";

cyclonev_ram_block ram_block1a16(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk0_output_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "rom";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "clock0";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 8191;
defparam ram_block1a16.port_a_logical_ram_depth = 65536;
defparam ram_block1a16.port_a_logical_ram_width = 24;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init3 = "000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a16.mem_init2 = "FFE000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFE00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFE00000000000000000000007FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFFFFFFFFFF80000000000000000000003FFFFFFFFFFFFFFFFFFFFFC";
defparam ram_block1a16.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFC0000000000000000000007FFFFFFFFFFFFFFFFFFFFF0000000000000000000001FFFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFFE000000000000000000000FFFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFF8000000000000000000003FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFFE000000000000000000003FFFFFFFFFFFFFFFFFFFF8";
defparam ram_block1a16.mem_init0 = "00000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000000";

cyclonev_ram_block ram_block1a40(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a40_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a40.clk0_core_clock_enable = "ena0";
defparam ram_block1a40.clk0_input_clock_enable = "ena0";
defparam ram_block1a40.clk0_output_clock_enable = "ena0";
defparam ram_block1a40.data_interleave_offset_in_bits = 1;
defparam ram_block1a40.data_interleave_width_in_bits = 1;
defparam ram_block1a40.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a40.init_file_layout = "port_a";
defparam ram_block1a40.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a40.operation_mode = "rom";
defparam ram_block1a40.port_a_address_clear = "none";
defparam ram_block1a40.port_a_address_width = 13;
defparam ram_block1a40.port_a_data_out_clear = "none";
defparam ram_block1a40.port_a_data_out_clock = "clock0";
defparam ram_block1a40.port_a_data_width = 1;
defparam ram_block1a40.port_a_first_address = 8192;
defparam ram_block1a40.port_a_first_bit_number = 16;
defparam ram_block1a40.port_a_last_address = 16383;
defparam ram_block1a40.port_a_logical_ram_depth = 65536;
defparam ram_block1a40.port_a_logical_ram_width = 24;
defparam ram_block1a40.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a40.ram_block_type = "auto";
defparam ram_block1a40.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a40.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000";
defparam ram_block1a40.mem_init1 = "00000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000";
defparam ram_block1a40.mem_init0 = "0000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000";

cyclonev_ram_block ram_block1a113(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a113_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a113.clk0_core_clock_enable = "ena0";
defparam ram_block1a113.clk0_input_clock_enable = "ena0";
defparam ram_block1a113.clk0_output_clock_enable = "ena0";
defparam ram_block1a113.data_interleave_offset_in_bits = 1;
defparam ram_block1a113.data_interleave_width_in_bits = 1;
defparam ram_block1a113.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a113.init_file_layout = "port_a";
defparam ram_block1a113.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a113.operation_mode = "rom";
defparam ram_block1a113.port_a_address_clear = "none";
defparam ram_block1a113.port_a_address_width = 13;
defparam ram_block1a113.port_a_data_out_clear = "none";
defparam ram_block1a113.port_a_data_out_clock = "clock0";
defparam ram_block1a113.port_a_data_width = 1;
defparam ram_block1a113.port_a_first_address = 32768;
defparam ram_block1a113.port_a_first_bit_number = 17;
defparam ram_block1a113.port_a_last_address = 40959;
defparam ram_block1a113.port_a_logical_ram_depth = 65536;
defparam ram_block1a113.port_a_logical_ram_width = 24;
defparam ram_block1a113.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a113.ram_block_type = "auto";
defparam ram_block1a113.mem_init3 = "000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000";
defparam ram_block1a113.mem_init2 = "000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a113.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a113.mem_init0 = "FFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

cyclonev_ram_block ram_block1a137(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a137_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a137.clk0_core_clock_enable = "ena0";
defparam ram_block1a137.clk0_input_clock_enable = "ena0";
defparam ram_block1a137.clk0_output_clock_enable = "ena0";
defparam ram_block1a137.data_interleave_offset_in_bits = 1;
defparam ram_block1a137.data_interleave_width_in_bits = 1;
defparam ram_block1a137.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a137.init_file_layout = "port_a";
defparam ram_block1a137.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a137.operation_mode = "rom";
defparam ram_block1a137.port_a_address_clear = "none";
defparam ram_block1a137.port_a_address_width = 13;
defparam ram_block1a137.port_a_data_out_clear = "none";
defparam ram_block1a137.port_a_data_out_clock = "clock0";
defparam ram_block1a137.port_a_data_width = 1;
defparam ram_block1a137.port_a_first_address = 40960;
defparam ram_block1a137.port_a_first_bit_number = 17;
defparam ram_block1a137.port_a_last_address = 49151;
defparam ram_block1a137.port_a_logical_ram_depth = 65536;
defparam ram_block1a137.port_a_logical_ram_width = 24;
defparam ram_block1a137.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a137.ram_block_type = "auto";
defparam ram_block1a137.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a137.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a137.mem_init1 = "00000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a137.mem_init0 = "0000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a161(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a161_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a161.clk0_core_clock_enable = "ena0";
defparam ram_block1a161.clk0_input_clock_enable = "ena0";
defparam ram_block1a161.clk0_output_clock_enable = "ena0";
defparam ram_block1a161.data_interleave_offset_in_bits = 1;
defparam ram_block1a161.data_interleave_width_in_bits = 1;
defparam ram_block1a161.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a161.init_file_layout = "port_a";
defparam ram_block1a161.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a161.operation_mode = "rom";
defparam ram_block1a161.port_a_address_clear = "none";
defparam ram_block1a161.port_a_address_width = 13;
defparam ram_block1a161.port_a_data_out_clear = "none";
defparam ram_block1a161.port_a_data_out_clock = "clock0";
defparam ram_block1a161.port_a_data_width = 1;
defparam ram_block1a161.port_a_first_address = 49152;
defparam ram_block1a161.port_a_first_bit_number = 17;
defparam ram_block1a161.port_a_last_address = 57343;
defparam ram_block1a161.port_a_logical_ram_depth = 65536;
defparam ram_block1a161.port_a_logical_ram_width = 24;
defparam ram_block1a161.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a161.ram_block_type = "auto";
defparam ram_block1a161.mem_init3 = "00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000";
defparam ram_block1a161.mem_init2 = "00000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000";
defparam ram_block1a161.mem_init1 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a161.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a185(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a185_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a185.clk0_core_clock_enable = "ena0";
defparam ram_block1a185.clk0_input_clock_enable = "ena0";
defparam ram_block1a185.clk0_output_clock_enable = "ena0";
defparam ram_block1a185.data_interleave_offset_in_bits = 1;
defparam ram_block1a185.data_interleave_width_in_bits = 1;
defparam ram_block1a185.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a185.init_file_layout = "port_a";
defparam ram_block1a185.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a185.operation_mode = "rom";
defparam ram_block1a185.port_a_address_clear = "none";
defparam ram_block1a185.port_a_address_width = 13;
defparam ram_block1a185.port_a_data_out_clear = "none";
defparam ram_block1a185.port_a_data_out_clock = "clock0";
defparam ram_block1a185.port_a_data_width = 1;
defparam ram_block1a185.port_a_first_address = 57344;
defparam ram_block1a185.port_a_first_bit_number = 17;
defparam ram_block1a185.port_a_last_address = 65535;
defparam ram_block1a185.port_a_logical_ram_depth = 65536;
defparam ram_block1a185.port_a_logical_ram_width = 24;
defparam ram_block1a185.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a185.ram_block_type = "auto";
defparam ram_block1a185.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a185.mem_init2 = "FFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a185.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000";
defparam ram_block1a185.mem_init0 = "0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000";

cyclonev_ram_block ram_block1a65(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a65_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a65.clk0_core_clock_enable = "ena0";
defparam ram_block1a65.clk0_input_clock_enable = "ena0";
defparam ram_block1a65.clk0_output_clock_enable = "ena0";
defparam ram_block1a65.data_interleave_offset_in_bits = 1;
defparam ram_block1a65.data_interleave_width_in_bits = 1;
defparam ram_block1a65.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a65.init_file_layout = "port_a";
defparam ram_block1a65.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a65.operation_mode = "rom";
defparam ram_block1a65.port_a_address_clear = "none";
defparam ram_block1a65.port_a_address_width = 13;
defparam ram_block1a65.port_a_data_out_clear = "none";
defparam ram_block1a65.port_a_data_out_clock = "clock0";
defparam ram_block1a65.port_a_data_width = 1;
defparam ram_block1a65.port_a_first_address = 16384;
defparam ram_block1a65.port_a_first_bit_number = 17;
defparam ram_block1a65.port_a_last_address = 24575;
defparam ram_block1a65.port_a_logical_ram_depth = 65536;
defparam ram_block1a65.port_a_logical_ram_width = 24;
defparam ram_block1a65.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a65.ram_block_type = "auto";
defparam ram_block1a65.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFF";
defparam ram_block1a65.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFF";
defparam ram_block1a65.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a65.mem_init0 = "000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a89(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a89_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a89.clk0_core_clock_enable = "ena0";
defparam ram_block1a89.clk0_input_clock_enable = "ena0";
defparam ram_block1a89.clk0_output_clock_enable = "ena0";
defparam ram_block1a89.data_interleave_offset_in_bits = 1;
defparam ram_block1a89.data_interleave_width_in_bits = 1;
defparam ram_block1a89.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a89.init_file_layout = "port_a";
defparam ram_block1a89.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a89.operation_mode = "rom";
defparam ram_block1a89.port_a_address_clear = "none";
defparam ram_block1a89.port_a_address_width = 13;
defparam ram_block1a89.port_a_data_out_clear = "none";
defparam ram_block1a89.port_a_data_out_clock = "clock0";
defparam ram_block1a89.port_a_data_width = 1;
defparam ram_block1a89.port_a_first_address = 24576;
defparam ram_block1a89.port_a_first_bit_number = 17;
defparam ram_block1a89.port_a_last_address = 32767;
defparam ram_block1a89.port_a_logical_ram_depth = 65536;
defparam ram_block1a89.port_a_logical_ram_width = 24;
defparam ram_block1a89.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a89.ram_block_type = "auto";
defparam ram_block1a89.mem_init3 = "00000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000";
defparam ram_block1a89.mem_init2 = "0000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a89.mem_init1 = "00000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a89.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a17(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk0_output_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "rom";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "clock0";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 8191;
defparam ram_block1a17.port_a_logical_ram_depth = 65536;
defparam ram_block1a17.port_a_logical_ram_width = 24;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init3 = "FFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a17.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000";
defparam ram_block1a17.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000";
defparam ram_block1a17.mem_init0 = "00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a41(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a41_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a41.clk0_core_clock_enable = "ena0";
defparam ram_block1a41.clk0_input_clock_enable = "ena0";
defparam ram_block1a41.clk0_output_clock_enable = "ena0";
defparam ram_block1a41.data_interleave_offset_in_bits = 1;
defparam ram_block1a41.data_interleave_width_in_bits = 1;
defparam ram_block1a41.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a41.init_file_layout = "port_a";
defparam ram_block1a41.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a41.operation_mode = "rom";
defparam ram_block1a41.port_a_address_clear = "none";
defparam ram_block1a41.port_a_address_width = 13;
defparam ram_block1a41.port_a_data_out_clear = "none";
defparam ram_block1a41.port_a_data_out_clock = "clock0";
defparam ram_block1a41.port_a_data_width = 1;
defparam ram_block1a41.port_a_first_address = 8192;
defparam ram_block1a41.port_a_first_bit_number = 17;
defparam ram_block1a41.port_a_last_address = 16383;
defparam ram_block1a41.port_a_logical_ram_depth = 65536;
defparam ram_block1a41.port_a_logical_ram_width = 24;
defparam ram_block1a41.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a41.ram_block_type = "auto";
defparam ram_block1a41.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000";
defparam ram_block1a41.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a41.mem_init1 = "FFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a41.mem_init0 = "FFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a114(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a114_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a114.clk0_core_clock_enable = "ena0";
defparam ram_block1a114.clk0_input_clock_enable = "ena0";
defparam ram_block1a114.clk0_output_clock_enable = "ena0";
defparam ram_block1a114.data_interleave_offset_in_bits = 1;
defparam ram_block1a114.data_interleave_width_in_bits = 1;
defparam ram_block1a114.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a114.init_file_layout = "port_a";
defparam ram_block1a114.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a114.operation_mode = "rom";
defparam ram_block1a114.port_a_address_clear = "none";
defparam ram_block1a114.port_a_address_width = 13;
defparam ram_block1a114.port_a_data_out_clear = "none";
defparam ram_block1a114.port_a_data_out_clock = "clock0";
defparam ram_block1a114.port_a_data_width = 1;
defparam ram_block1a114.port_a_first_address = 32768;
defparam ram_block1a114.port_a_first_bit_number = 18;
defparam ram_block1a114.port_a_last_address = 40959;
defparam ram_block1a114.port_a_logical_ram_depth = 65536;
defparam ram_block1a114.port_a_logical_ram_width = 24;
defparam ram_block1a114.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a114.ram_block_type = "auto";
defparam ram_block1a114.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000";
defparam ram_block1a114.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a114.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a114.mem_init0 = "FFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

cyclonev_ram_block ram_block1a138(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a138_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a138.clk0_core_clock_enable = "ena0";
defparam ram_block1a138.clk0_input_clock_enable = "ena0";
defparam ram_block1a138.clk0_output_clock_enable = "ena0";
defparam ram_block1a138.data_interleave_offset_in_bits = 1;
defparam ram_block1a138.data_interleave_width_in_bits = 1;
defparam ram_block1a138.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a138.init_file_layout = "port_a";
defparam ram_block1a138.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a138.operation_mode = "rom";
defparam ram_block1a138.port_a_address_clear = "none";
defparam ram_block1a138.port_a_address_width = 13;
defparam ram_block1a138.port_a_data_out_clear = "none";
defparam ram_block1a138.port_a_data_out_clock = "clock0";
defparam ram_block1a138.port_a_data_width = 1;
defparam ram_block1a138.port_a_first_address = 40960;
defparam ram_block1a138.port_a_first_bit_number = 18;
defparam ram_block1a138.port_a_last_address = 49151;
defparam ram_block1a138.port_a_logical_ram_depth = 65536;
defparam ram_block1a138.port_a_logical_ram_width = 24;
defparam ram_block1a138.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a138.ram_block_type = "auto";
defparam ram_block1a138.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a138.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a138.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a138.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a162(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a162_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a162.clk0_core_clock_enable = "ena0";
defparam ram_block1a162.clk0_input_clock_enable = "ena0";
defparam ram_block1a162.clk0_output_clock_enable = "ena0";
defparam ram_block1a162.data_interleave_offset_in_bits = 1;
defparam ram_block1a162.data_interleave_width_in_bits = 1;
defparam ram_block1a162.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a162.init_file_layout = "port_a";
defparam ram_block1a162.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a162.operation_mode = "rom";
defparam ram_block1a162.port_a_address_clear = "none";
defparam ram_block1a162.port_a_address_width = 13;
defparam ram_block1a162.port_a_data_out_clear = "none";
defparam ram_block1a162.port_a_data_out_clock = "clock0";
defparam ram_block1a162.port_a_data_width = 1;
defparam ram_block1a162.port_a_first_address = 49152;
defparam ram_block1a162.port_a_first_bit_number = 18;
defparam ram_block1a162.port_a_last_address = 57343;
defparam ram_block1a162.port_a_logical_ram_depth = 65536;
defparam ram_block1a162.port_a_logical_ram_width = 24;
defparam ram_block1a162.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a162.ram_block_type = "auto";
defparam ram_block1a162.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a162.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a162.mem_init1 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a162.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a186(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a186_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a186.clk0_core_clock_enable = "ena0";
defparam ram_block1a186.clk0_input_clock_enable = "ena0";
defparam ram_block1a186.clk0_output_clock_enable = "ena0";
defparam ram_block1a186.data_interleave_offset_in_bits = 1;
defparam ram_block1a186.data_interleave_width_in_bits = 1;
defparam ram_block1a186.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a186.init_file_layout = "port_a";
defparam ram_block1a186.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a186.operation_mode = "rom";
defparam ram_block1a186.port_a_address_clear = "none";
defparam ram_block1a186.port_a_address_width = 13;
defparam ram_block1a186.port_a_data_out_clear = "none";
defparam ram_block1a186.port_a_data_out_clock = "clock0";
defparam ram_block1a186.port_a_data_width = 1;
defparam ram_block1a186.port_a_first_address = 57344;
defparam ram_block1a186.port_a_first_bit_number = 18;
defparam ram_block1a186.port_a_last_address = 65535;
defparam ram_block1a186.port_a_logical_ram_depth = 65536;
defparam ram_block1a186.port_a_logical_ram_width = 24;
defparam ram_block1a186.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a186.ram_block_type = "auto";
defparam ram_block1a186.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a186.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a186.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a186.mem_init0 = "0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a66(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a66_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a66.clk0_core_clock_enable = "ena0";
defparam ram_block1a66.clk0_input_clock_enable = "ena0";
defparam ram_block1a66.clk0_output_clock_enable = "ena0";
defparam ram_block1a66.data_interleave_offset_in_bits = 1;
defparam ram_block1a66.data_interleave_width_in_bits = 1;
defparam ram_block1a66.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a66.init_file_layout = "port_a";
defparam ram_block1a66.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a66.operation_mode = "rom";
defparam ram_block1a66.port_a_address_clear = "none";
defparam ram_block1a66.port_a_address_width = 13;
defparam ram_block1a66.port_a_data_out_clear = "none";
defparam ram_block1a66.port_a_data_out_clock = "clock0";
defparam ram_block1a66.port_a_data_width = 1;
defparam ram_block1a66.port_a_first_address = 16384;
defparam ram_block1a66.port_a_first_bit_number = 18;
defparam ram_block1a66.port_a_last_address = 24575;
defparam ram_block1a66.port_a_logical_ram_depth = 65536;
defparam ram_block1a66.port_a_logical_ram_width = 24;
defparam ram_block1a66.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a66.ram_block_type = "auto";
defparam ram_block1a66.mem_init3 = "00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a66.mem_init2 = "00000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a66.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a66.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a90(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a90_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a90.clk0_core_clock_enable = "ena0";
defparam ram_block1a90.clk0_input_clock_enable = "ena0";
defparam ram_block1a90.clk0_output_clock_enable = "ena0";
defparam ram_block1a90.data_interleave_offset_in_bits = 1;
defparam ram_block1a90.data_interleave_width_in_bits = 1;
defparam ram_block1a90.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a90.init_file_layout = "port_a";
defparam ram_block1a90.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a90.operation_mode = "rom";
defparam ram_block1a90.port_a_address_clear = "none";
defparam ram_block1a90.port_a_address_width = 13;
defparam ram_block1a90.port_a_data_out_clear = "none";
defparam ram_block1a90.port_a_data_out_clock = "clock0";
defparam ram_block1a90.port_a_data_width = 1;
defparam ram_block1a90.port_a_first_address = 24576;
defparam ram_block1a90.port_a_first_bit_number = 18;
defparam ram_block1a90.port_a_last_address = 32767;
defparam ram_block1a90.port_a_logical_ram_depth = 65536;
defparam ram_block1a90.port_a_logical_ram_width = 24;
defparam ram_block1a90.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a90.ram_block_type = "auto";
defparam ram_block1a90.mem_init3 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000";
defparam ram_block1a90.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a90.mem_init1 = "0000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a90.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a18(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk0_output_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "rom";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "clock0";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 8191;
defparam ram_block1a18.port_a_logical_ram_depth = 65536;
defparam ram_block1a18.port_a_logical_ram_width = 24;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a18.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init0 = "00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a42(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a42_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a42.clk0_core_clock_enable = "ena0";
defparam ram_block1a42.clk0_input_clock_enable = "ena0";
defparam ram_block1a42.clk0_output_clock_enable = "ena0";
defparam ram_block1a42.data_interleave_offset_in_bits = 1;
defparam ram_block1a42.data_interleave_width_in_bits = 1;
defparam ram_block1a42.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a42.init_file_layout = "port_a";
defparam ram_block1a42.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a42.operation_mode = "rom";
defparam ram_block1a42.port_a_address_clear = "none";
defparam ram_block1a42.port_a_address_width = 13;
defparam ram_block1a42.port_a_data_out_clear = "none";
defparam ram_block1a42.port_a_data_out_clock = "clock0";
defparam ram_block1a42.port_a_data_width = 1;
defparam ram_block1a42.port_a_first_address = 8192;
defparam ram_block1a42.port_a_first_bit_number = 18;
defparam ram_block1a42.port_a_last_address = 16383;
defparam ram_block1a42.port_a_logical_ram_depth = 65536;
defparam ram_block1a42.port_a_logical_ram_width = 24;
defparam ram_block1a42.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a42.ram_block_type = "auto";
defparam ram_block1a42.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a42.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a42.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a42.mem_init0 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a115(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a115_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a115.clk0_core_clock_enable = "ena0";
defparam ram_block1a115.clk0_input_clock_enable = "ena0";
defparam ram_block1a115.clk0_output_clock_enable = "ena0";
defparam ram_block1a115.data_interleave_offset_in_bits = 1;
defparam ram_block1a115.data_interleave_width_in_bits = 1;
defparam ram_block1a115.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a115.init_file_layout = "port_a";
defparam ram_block1a115.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a115.operation_mode = "rom";
defparam ram_block1a115.port_a_address_clear = "none";
defparam ram_block1a115.port_a_address_width = 13;
defparam ram_block1a115.port_a_data_out_clear = "none";
defparam ram_block1a115.port_a_data_out_clock = "clock0";
defparam ram_block1a115.port_a_data_width = 1;
defparam ram_block1a115.port_a_first_address = 32768;
defparam ram_block1a115.port_a_first_bit_number = 19;
defparam ram_block1a115.port_a_last_address = 40959;
defparam ram_block1a115.port_a_logical_ram_depth = 65536;
defparam ram_block1a115.port_a_logical_ram_width = 24;
defparam ram_block1a115.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a115.ram_block_type = "auto";
defparam ram_block1a115.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a115.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a115.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a115.mem_init0 = "00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

cyclonev_ram_block ram_block1a139(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a139_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a139.clk0_core_clock_enable = "ena0";
defparam ram_block1a139.clk0_input_clock_enable = "ena0";
defparam ram_block1a139.clk0_output_clock_enable = "ena0";
defparam ram_block1a139.data_interleave_offset_in_bits = 1;
defparam ram_block1a139.data_interleave_width_in_bits = 1;
defparam ram_block1a139.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a139.init_file_layout = "port_a";
defparam ram_block1a139.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a139.operation_mode = "rom";
defparam ram_block1a139.port_a_address_clear = "none";
defparam ram_block1a139.port_a_address_width = 13;
defparam ram_block1a139.port_a_data_out_clear = "none";
defparam ram_block1a139.port_a_data_out_clock = "clock0";
defparam ram_block1a139.port_a_data_width = 1;
defparam ram_block1a139.port_a_first_address = 40960;
defparam ram_block1a139.port_a_first_bit_number = 19;
defparam ram_block1a139.port_a_last_address = 49151;
defparam ram_block1a139.port_a_logical_ram_depth = 65536;
defparam ram_block1a139.port_a_logical_ram_width = 24;
defparam ram_block1a139.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a139.ram_block_type = "auto";
defparam ram_block1a139.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a139.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a139.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a139.mem_init0 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a163(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a163_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a163.clk0_core_clock_enable = "ena0";
defparam ram_block1a163.clk0_input_clock_enable = "ena0";
defparam ram_block1a163.clk0_output_clock_enable = "ena0";
defparam ram_block1a163.data_interleave_offset_in_bits = 1;
defparam ram_block1a163.data_interleave_width_in_bits = 1;
defparam ram_block1a163.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a163.init_file_layout = "port_a";
defparam ram_block1a163.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a163.operation_mode = "rom";
defparam ram_block1a163.port_a_address_clear = "none";
defparam ram_block1a163.port_a_address_width = 13;
defparam ram_block1a163.port_a_data_out_clear = "none";
defparam ram_block1a163.port_a_data_out_clock = "clock0";
defparam ram_block1a163.port_a_data_width = 1;
defparam ram_block1a163.port_a_first_address = 49152;
defparam ram_block1a163.port_a_first_bit_number = 19;
defparam ram_block1a163.port_a_last_address = 57343;
defparam ram_block1a163.port_a_logical_ram_depth = 65536;
defparam ram_block1a163.port_a_logical_ram_width = 24;
defparam ram_block1a163.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a163.ram_block_type = "auto";
defparam ram_block1a163.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a163.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a163.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a163.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a187(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a187_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a187.clk0_core_clock_enable = "ena0";
defparam ram_block1a187.clk0_input_clock_enable = "ena0";
defparam ram_block1a187.clk0_output_clock_enable = "ena0";
defparam ram_block1a187.data_interleave_offset_in_bits = 1;
defparam ram_block1a187.data_interleave_width_in_bits = 1;
defparam ram_block1a187.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a187.init_file_layout = "port_a";
defparam ram_block1a187.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a187.operation_mode = "rom";
defparam ram_block1a187.port_a_address_clear = "none";
defparam ram_block1a187.port_a_address_width = 13;
defparam ram_block1a187.port_a_data_out_clear = "none";
defparam ram_block1a187.port_a_data_out_clock = "clock0";
defparam ram_block1a187.port_a_data_width = 1;
defparam ram_block1a187.port_a_first_address = 57344;
defparam ram_block1a187.port_a_first_bit_number = 19;
defparam ram_block1a187.port_a_last_address = 65535;
defparam ram_block1a187.port_a_logical_ram_depth = 65536;
defparam ram_block1a187.port_a_logical_ram_width = 24;
defparam ram_block1a187.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a187.ram_block_type = "auto";
defparam ram_block1a187.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000";
defparam ram_block1a187.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a187.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a187.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a67(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a67_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a67.clk0_core_clock_enable = "ena0";
defparam ram_block1a67.clk0_input_clock_enable = "ena0";
defparam ram_block1a67.clk0_output_clock_enable = "ena0";
defparam ram_block1a67.data_interleave_offset_in_bits = 1;
defparam ram_block1a67.data_interleave_width_in_bits = 1;
defparam ram_block1a67.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a67.init_file_layout = "port_a";
defparam ram_block1a67.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a67.operation_mode = "rom";
defparam ram_block1a67.port_a_address_clear = "none";
defparam ram_block1a67.port_a_address_width = 13;
defparam ram_block1a67.port_a_data_out_clear = "none";
defparam ram_block1a67.port_a_data_out_clock = "clock0";
defparam ram_block1a67.port_a_data_width = 1;
defparam ram_block1a67.port_a_first_address = 16384;
defparam ram_block1a67.port_a_first_bit_number = 19;
defparam ram_block1a67.port_a_last_address = 24575;
defparam ram_block1a67.port_a_logical_ram_depth = 65536;
defparam ram_block1a67.port_a_logical_ram_width = 24;
defparam ram_block1a67.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a67.ram_block_type = "auto";
defparam ram_block1a67.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a67.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a67.mem_init1 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a67.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a91(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a91_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a91.clk0_core_clock_enable = "ena0";
defparam ram_block1a91.clk0_input_clock_enable = "ena0";
defparam ram_block1a91.clk0_output_clock_enable = "ena0";
defparam ram_block1a91.data_interleave_offset_in_bits = 1;
defparam ram_block1a91.data_interleave_width_in_bits = 1;
defparam ram_block1a91.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a91.init_file_layout = "port_a";
defparam ram_block1a91.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a91.operation_mode = "rom";
defparam ram_block1a91.port_a_address_clear = "none";
defparam ram_block1a91.port_a_address_width = 13;
defparam ram_block1a91.port_a_data_out_clear = "none";
defparam ram_block1a91.port_a_data_out_clock = "clock0";
defparam ram_block1a91.port_a_data_width = 1;
defparam ram_block1a91.port_a_first_address = 24576;
defparam ram_block1a91.port_a_first_bit_number = 19;
defparam ram_block1a91.port_a_last_address = 32767;
defparam ram_block1a91.port_a_logical_ram_depth = 65536;
defparam ram_block1a91.port_a_logical_ram_width = 24;
defparam ram_block1a91.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a91.ram_block_type = "auto";
defparam ram_block1a91.mem_init3 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a91.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a91.mem_init1 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a91.mem_init0 = "0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a19(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk0_output_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "rom";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "clock0";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 8191;
defparam ram_block1a19.port_a_logical_ram_depth = 65536;
defparam ram_block1a19.port_a_logical_ram_width = 24;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000";
defparam ram_block1a19.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a19.mem_init0 = "FFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a43(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a43_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a43.clk0_core_clock_enable = "ena0";
defparam ram_block1a43.clk0_input_clock_enable = "ena0";
defparam ram_block1a43.clk0_output_clock_enable = "ena0";
defparam ram_block1a43.data_interleave_offset_in_bits = 1;
defparam ram_block1a43.data_interleave_width_in_bits = 1;
defparam ram_block1a43.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a43.init_file_layout = "port_a";
defparam ram_block1a43.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a43.operation_mode = "rom";
defparam ram_block1a43.port_a_address_clear = "none";
defparam ram_block1a43.port_a_address_width = 13;
defparam ram_block1a43.port_a_data_out_clear = "none";
defparam ram_block1a43.port_a_data_out_clock = "clock0";
defparam ram_block1a43.port_a_data_width = 1;
defparam ram_block1a43.port_a_first_address = 8192;
defparam ram_block1a43.port_a_first_bit_number = 19;
defparam ram_block1a43.port_a_last_address = 16383;
defparam ram_block1a43.port_a_logical_ram_depth = 65536;
defparam ram_block1a43.port_a_logical_ram_width = 24;
defparam ram_block1a43.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a43.ram_block_type = "auto";
defparam ram_block1a43.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a43.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a43.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a43.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a116(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a116_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a116.clk0_core_clock_enable = "ena0";
defparam ram_block1a116.clk0_input_clock_enable = "ena0";
defparam ram_block1a116.clk0_output_clock_enable = "ena0";
defparam ram_block1a116.data_interleave_offset_in_bits = 1;
defparam ram_block1a116.data_interleave_width_in_bits = 1;
defparam ram_block1a116.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a116.init_file_layout = "port_a";
defparam ram_block1a116.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a116.operation_mode = "rom";
defparam ram_block1a116.port_a_address_clear = "none";
defparam ram_block1a116.port_a_address_width = 13;
defparam ram_block1a116.port_a_data_out_clear = "none";
defparam ram_block1a116.port_a_data_out_clock = "clock0";
defparam ram_block1a116.port_a_data_width = 1;
defparam ram_block1a116.port_a_first_address = 32768;
defparam ram_block1a116.port_a_first_bit_number = 20;
defparam ram_block1a116.port_a_last_address = 40959;
defparam ram_block1a116.port_a_logical_ram_depth = 65536;
defparam ram_block1a116.port_a_logical_ram_width = 24;
defparam ram_block1a116.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a116.ram_block_type = "auto";
defparam ram_block1a116.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a116.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a116.mem_init1 = "0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a116.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

cyclonev_ram_block ram_block1a140(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a140_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a140.clk0_core_clock_enable = "ena0";
defparam ram_block1a140.clk0_input_clock_enable = "ena0";
defparam ram_block1a140.clk0_output_clock_enable = "ena0";
defparam ram_block1a140.data_interleave_offset_in_bits = 1;
defparam ram_block1a140.data_interleave_width_in_bits = 1;
defparam ram_block1a140.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a140.init_file_layout = "port_a";
defparam ram_block1a140.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a140.operation_mode = "rom";
defparam ram_block1a140.port_a_address_clear = "none";
defparam ram_block1a140.port_a_address_width = 13;
defparam ram_block1a140.port_a_data_out_clear = "none";
defparam ram_block1a140.port_a_data_out_clock = "clock0";
defparam ram_block1a140.port_a_data_width = 1;
defparam ram_block1a140.port_a_first_address = 40960;
defparam ram_block1a140.port_a_first_bit_number = 20;
defparam ram_block1a140.port_a_last_address = 49151;
defparam ram_block1a140.port_a_logical_ram_depth = 65536;
defparam ram_block1a140.port_a_logical_ram_width = 24;
defparam ram_block1a140.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a140.ram_block_type = "auto";
defparam ram_block1a140.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a140.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a140.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a140.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a164(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a164_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a164.clk0_core_clock_enable = "ena0";
defparam ram_block1a164.clk0_input_clock_enable = "ena0";
defparam ram_block1a164.clk0_output_clock_enable = "ena0";
defparam ram_block1a164.data_interleave_offset_in_bits = 1;
defparam ram_block1a164.data_interleave_width_in_bits = 1;
defparam ram_block1a164.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a164.init_file_layout = "port_a";
defparam ram_block1a164.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a164.operation_mode = "rom";
defparam ram_block1a164.port_a_address_clear = "none";
defparam ram_block1a164.port_a_address_width = 13;
defparam ram_block1a164.port_a_data_out_clear = "none";
defparam ram_block1a164.port_a_data_out_clock = "clock0";
defparam ram_block1a164.port_a_data_width = 1;
defparam ram_block1a164.port_a_first_address = 49152;
defparam ram_block1a164.port_a_first_bit_number = 20;
defparam ram_block1a164.port_a_last_address = 57343;
defparam ram_block1a164.port_a_logical_ram_depth = 65536;
defparam ram_block1a164.port_a_logical_ram_width = 24;
defparam ram_block1a164.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a164.ram_block_type = "auto";
defparam ram_block1a164.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a164.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a164.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a164.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a188(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a188_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a188.clk0_core_clock_enable = "ena0";
defparam ram_block1a188.clk0_input_clock_enable = "ena0";
defparam ram_block1a188.clk0_output_clock_enable = "ena0";
defparam ram_block1a188.data_interleave_offset_in_bits = 1;
defparam ram_block1a188.data_interleave_width_in_bits = 1;
defparam ram_block1a188.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a188.init_file_layout = "port_a";
defparam ram_block1a188.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a188.operation_mode = "rom";
defparam ram_block1a188.port_a_address_clear = "none";
defparam ram_block1a188.port_a_address_width = 13;
defparam ram_block1a188.port_a_data_out_clear = "none";
defparam ram_block1a188.port_a_data_out_clock = "clock0";
defparam ram_block1a188.port_a_data_width = 1;
defparam ram_block1a188.port_a_first_address = 57344;
defparam ram_block1a188.port_a_first_bit_number = 20;
defparam ram_block1a188.port_a_last_address = 65535;
defparam ram_block1a188.port_a_logical_ram_depth = 65536;
defparam ram_block1a188.port_a_logical_ram_width = 24;
defparam ram_block1a188.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a188.ram_block_type = "auto";
defparam ram_block1a188.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a188.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000";
defparam ram_block1a188.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a188.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a68(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a68_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a68.clk0_core_clock_enable = "ena0";
defparam ram_block1a68.clk0_input_clock_enable = "ena0";
defparam ram_block1a68.clk0_output_clock_enable = "ena0";
defparam ram_block1a68.data_interleave_offset_in_bits = 1;
defparam ram_block1a68.data_interleave_width_in_bits = 1;
defparam ram_block1a68.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a68.init_file_layout = "port_a";
defparam ram_block1a68.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a68.operation_mode = "rom";
defparam ram_block1a68.port_a_address_clear = "none";
defparam ram_block1a68.port_a_address_width = 13;
defparam ram_block1a68.port_a_data_out_clear = "none";
defparam ram_block1a68.port_a_data_out_clock = "clock0";
defparam ram_block1a68.port_a_data_width = 1;
defparam ram_block1a68.port_a_first_address = 16384;
defparam ram_block1a68.port_a_first_bit_number = 20;
defparam ram_block1a68.port_a_last_address = 24575;
defparam ram_block1a68.port_a_logical_ram_depth = 65536;
defparam ram_block1a68.port_a_logical_ram_width = 24;
defparam ram_block1a68.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a68.ram_block_type = "auto";
defparam ram_block1a68.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a68.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a68.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a68.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a92(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a92_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a92.clk0_core_clock_enable = "ena0";
defparam ram_block1a92.clk0_input_clock_enable = "ena0";
defparam ram_block1a92.clk0_output_clock_enable = "ena0";
defparam ram_block1a92.data_interleave_offset_in_bits = 1;
defparam ram_block1a92.data_interleave_width_in_bits = 1;
defparam ram_block1a92.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a92.init_file_layout = "port_a";
defparam ram_block1a92.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a92.operation_mode = "rom";
defparam ram_block1a92.port_a_address_clear = "none";
defparam ram_block1a92.port_a_address_width = 13;
defparam ram_block1a92.port_a_data_out_clear = "none";
defparam ram_block1a92.port_a_data_out_clock = "clock0";
defparam ram_block1a92.port_a_data_width = 1;
defparam ram_block1a92.port_a_first_address = 24576;
defparam ram_block1a92.port_a_first_bit_number = 20;
defparam ram_block1a92.port_a_last_address = 32767;
defparam ram_block1a92.port_a_logical_ram_depth = 65536;
defparam ram_block1a92.port_a_logical_ram_width = 24;
defparam ram_block1a92.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a92.ram_block_type = "auto";
defparam ram_block1a92.mem_init3 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a92.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a92.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a92.mem_init0 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a20(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.clk0_output_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "rom";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "clock0";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 8191;
defparam ram_block1a20.port_a_logical_ram_depth = 65536;
defparam ram_block1a20.port_a_logical_ram_width = 24;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a20.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a20.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a44(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a44_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a44.clk0_core_clock_enable = "ena0";
defparam ram_block1a44.clk0_input_clock_enable = "ena0";
defparam ram_block1a44.clk0_output_clock_enable = "ena0";
defparam ram_block1a44.data_interleave_offset_in_bits = 1;
defparam ram_block1a44.data_interleave_width_in_bits = 1;
defparam ram_block1a44.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a44.init_file_layout = "port_a";
defparam ram_block1a44.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a44.operation_mode = "rom";
defparam ram_block1a44.port_a_address_clear = "none";
defparam ram_block1a44.port_a_address_width = 13;
defparam ram_block1a44.port_a_data_out_clear = "none";
defparam ram_block1a44.port_a_data_out_clock = "clock0";
defparam ram_block1a44.port_a_data_width = 1;
defparam ram_block1a44.port_a_first_address = 8192;
defparam ram_block1a44.port_a_first_bit_number = 20;
defparam ram_block1a44.port_a_last_address = 16383;
defparam ram_block1a44.port_a_logical_ram_depth = 65536;
defparam ram_block1a44.port_a_logical_ram_width = 24;
defparam ram_block1a44.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a44.ram_block_type = "auto";
defparam ram_block1a44.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a44.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a44.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a44.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a117(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a117_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a117.clk0_core_clock_enable = "ena0";
defparam ram_block1a117.clk0_input_clock_enable = "ena0";
defparam ram_block1a117.clk0_output_clock_enable = "ena0";
defparam ram_block1a117.data_interleave_offset_in_bits = 1;
defparam ram_block1a117.data_interleave_width_in_bits = 1;
defparam ram_block1a117.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a117.init_file_layout = "port_a";
defparam ram_block1a117.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a117.operation_mode = "rom";
defparam ram_block1a117.port_a_address_clear = "none";
defparam ram_block1a117.port_a_address_width = 13;
defparam ram_block1a117.port_a_data_out_clear = "none";
defparam ram_block1a117.port_a_data_out_clock = "clock0";
defparam ram_block1a117.port_a_data_width = 1;
defparam ram_block1a117.port_a_first_address = 32768;
defparam ram_block1a117.port_a_first_bit_number = 21;
defparam ram_block1a117.port_a_last_address = 40959;
defparam ram_block1a117.port_a_logical_ram_depth = 65536;
defparam ram_block1a117.port_a_logical_ram_width = 24;
defparam ram_block1a117.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a117.ram_block_type = "auto";
defparam ram_block1a117.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a117.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a117.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a117.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

cyclonev_ram_block ram_block1a141(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a141_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a141.clk0_core_clock_enable = "ena0";
defparam ram_block1a141.clk0_input_clock_enable = "ena0";
defparam ram_block1a141.clk0_output_clock_enable = "ena0";
defparam ram_block1a141.data_interleave_offset_in_bits = 1;
defparam ram_block1a141.data_interleave_width_in_bits = 1;
defparam ram_block1a141.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a141.init_file_layout = "port_a";
defparam ram_block1a141.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a141.operation_mode = "rom";
defparam ram_block1a141.port_a_address_clear = "none";
defparam ram_block1a141.port_a_address_width = 13;
defparam ram_block1a141.port_a_data_out_clear = "none";
defparam ram_block1a141.port_a_data_out_clock = "clock0";
defparam ram_block1a141.port_a_data_width = 1;
defparam ram_block1a141.port_a_first_address = 40960;
defparam ram_block1a141.port_a_first_bit_number = 21;
defparam ram_block1a141.port_a_last_address = 49151;
defparam ram_block1a141.port_a_logical_ram_depth = 65536;
defparam ram_block1a141.port_a_logical_ram_width = 24;
defparam ram_block1a141.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a141.ram_block_type = "auto";
defparam ram_block1a141.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a141.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a141.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a141.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a165(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a165_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a165.clk0_core_clock_enable = "ena0";
defparam ram_block1a165.clk0_input_clock_enable = "ena0";
defparam ram_block1a165.clk0_output_clock_enable = "ena0";
defparam ram_block1a165.data_interleave_offset_in_bits = 1;
defparam ram_block1a165.data_interleave_width_in_bits = 1;
defparam ram_block1a165.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a165.init_file_layout = "port_a";
defparam ram_block1a165.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a165.operation_mode = "rom";
defparam ram_block1a165.port_a_address_clear = "none";
defparam ram_block1a165.port_a_address_width = 13;
defparam ram_block1a165.port_a_data_out_clear = "none";
defparam ram_block1a165.port_a_data_out_clock = "clock0";
defparam ram_block1a165.port_a_data_width = 1;
defparam ram_block1a165.port_a_first_address = 49152;
defparam ram_block1a165.port_a_first_bit_number = 21;
defparam ram_block1a165.port_a_last_address = 57343;
defparam ram_block1a165.port_a_logical_ram_depth = 65536;
defparam ram_block1a165.port_a_logical_ram_width = 24;
defparam ram_block1a165.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a165.ram_block_type = "auto";
defparam ram_block1a165.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a165.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a165.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a165.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a189(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a189_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a189.clk0_core_clock_enable = "ena0";
defparam ram_block1a189.clk0_input_clock_enable = "ena0";
defparam ram_block1a189.clk0_output_clock_enable = "ena0";
defparam ram_block1a189.data_interleave_offset_in_bits = 1;
defparam ram_block1a189.data_interleave_width_in_bits = 1;
defparam ram_block1a189.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a189.init_file_layout = "port_a";
defparam ram_block1a189.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a189.operation_mode = "rom";
defparam ram_block1a189.port_a_address_clear = "none";
defparam ram_block1a189.port_a_address_width = 13;
defparam ram_block1a189.port_a_data_out_clear = "none";
defparam ram_block1a189.port_a_data_out_clock = "clock0";
defparam ram_block1a189.port_a_data_width = 1;
defparam ram_block1a189.port_a_first_address = 57344;
defparam ram_block1a189.port_a_first_bit_number = 21;
defparam ram_block1a189.port_a_last_address = 65535;
defparam ram_block1a189.port_a_logical_ram_depth = 65536;
defparam ram_block1a189.port_a_logical_ram_width = 24;
defparam ram_block1a189.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a189.ram_block_type = "auto";
defparam ram_block1a189.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a189.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a189.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a189.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a69(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a69_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a69.clk0_core_clock_enable = "ena0";
defparam ram_block1a69.clk0_input_clock_enable = "ena0";
defparam ram_block1a69.clk0_output_clock_enable = "ena0";
defparam ram_block1a69.data_interleave_offset_in_bits = 1;
defparam ram_block1a69.data_interleave_width_in_bits = 1;
defparam ram_block1a69.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a69.init_file_layout = "port_a";
defparam ram_block1a69.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a69.operation_mode = "rom";
defparam ram_block1a69.port_a_address_clear = "none";
defparam ram_block1a69.port_a_address_width = 13;
defparam ram_block1a69.port_a_data_out_clear = "none";
defparam ram_block1a69.port_a_data_out_clock = "clock0";
defparam ram_block1a69.port_a_data_width = 1;
defparam ram_block1a69.port_a_first_address = 16384;
defparam ram_block1a69.port_a_first_bit_number = 21;
defparam ram_block1a69.port_a_last_address = 24575;
defparam ram_block1a69.port_a_logical_ram_depth = 65536;
defparam ram_block1a69.port_a_logical_ram_width = 24;
defparam ram_block1a69.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a69.ram_block_type = "auto";
defparam ram_block1a69.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a69.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a69.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a69.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a93(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a93_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a93.clk0_core_clock_enable = "ena0";
defparam ram_block1a93.clk0_input_clock_enable = "ena0";
defparam ram_block1a93.clk0_output_clock_enable = "ena0";
defparam ram_block1a93.data_interleave_offset_in_bits = 1;
defparam ram_block1a93.data_interleave_width_in_bits = 1;
defparam ram_block1a93.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a93.init_file_layout = "port_a";
defparam ram_block1a93.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a93.operation_mode = "rom";
defparam ram_block1a93.port_a_address_clear = "none";
defparam ram_block1a93.port_a_address_width = 13;
defparam ram_block1a93.port_a_data_out_clear = "none";
defparam ram_block1a93.port_a_data_out_clock = "clock0";
defparam ram_block1a93.port_a_data_width = 1;
defparam ram_block1a93.port_a_first_address = 24576;
defparam ram_block1a93.port_a_first_bit_number = 21;
defparam ram_block1a93.port_a_last_address = 32767;
defparam ram_block1a93.port_a_logical_ram_depth = 65536;
defparam ram_block1a93.port_a_logical_ram_width = 24;
defparam ram_block1a93.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a93.ram_block_type = "auto";
defparam ram_block1a93.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a93.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a93.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a93.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a21(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.clk0_output_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "rom";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "clock0";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 8191;
defparam ram_block1a21.port_a_logical_ram_depth = 65536;
defparam ram_block1a21.port_a_logical_ram_width = 24;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a21.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a45(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a45_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a45.clk0_core_clock_enable = "ena0";
defparam ram_block1a45.clk0_input_clock_enable = "ena0";
defparam ram_block1a45.clk0_output_clock_enable = "ena0";
defparam ram_block1a45.data_interleave_offset_in_bits = 1;
defparam ram_block1a45.data_interleave_width_in_bits = 1;
defparam ram_block1a45.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a45.init_file_layout = "port_a";
defparam ram_block1a45.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a45.operation_mode = "rom";
defparam ram_block1a45.port_a_address_clear = "none";
defparam ram_block1a45.port_a_address_width = 13;
defparam ram_block1a45.port_a_data_out_clear = "none";
defparam ram_block1a45.port_a_data_out_clock = "clock0";
defparam ram_block1a45.port_a_data_width = 1;
defparam ram_block1a45.port_a_first_address = 8192;
defparam ram_block1a45.port_a_first_bit_number = 21;
defparam ram_block1a45.port_a_last_address = 16383;
defparam ram_block1a45.port_a_logical_ram_depth = 65536;
defparam ram_block1a45.port_a_logical_ram_width = 24;
defparam ram_block1a45.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a45.ram_block_type = "auto";
defparam ram_block1a45.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a45.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a45.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a45.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a118(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a118_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a118.clk0_core_clock_enable = "ena0";
defparam ram_block1a118.clk0_input_clock_enable = "ena0";
defparam ram_block1a118.clk0_output_clock_enable = "ena0";
defparam ram_block1a118.data_interleave_offset_in_bits = 1;
defparam ram_block1a118.data_interleave_width_in_bits = 1;
defparam ram_block1a118.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a118.init_file_layout = "port_a";
defparam ram_block1a118.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a118.operation_mode = "rom";
defparam ram_block1a118.port_a_address_clear = "none";
defparam ram_block1a118.port_a_address_width = 13;
defparam ram_block1a118.port_a_data_out_clear = "none";
defparam ram_block1a118.port_a_data_out_clock = "clock0";
defparam ram_block1a118.port_a_data_width = 1;
defparam ram_block1a118.port_a_first_address = 32768;
defparam ram_block1a118.port_a_first_bit_number = 22;
defparam ram_block1a118.port_a_last_address = 40959;
defparam ram_block1a118.port_a_logical_ram_depth = 65536;
defparam ram_block1a118.port_a_logical_ram_width = 24;
defparam ram_block1a118.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a118.ram_block_type = "auto";
defparam ram_block1a118.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a118.mem_init2 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a118.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a118.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

cyclonev_ram_block ram_block1a142(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a142_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a142.clk0_core_clock_enable = "ena0";
defparam ram_block1a142.clk0_input_clock_enable = "ena0";
defparam ram_block1a142.clk0_output_clock_enable = "ena0";
defparam ram_block1a142.data_interleave_offset_in_bits = 1;
defparam ram_block1a142.data_interleave_width_in_bits = 1;
defparam ram_block1a142.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a142.init_file_layout = "port_a";
defparam ram_block1a142.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a142.operation_mode = "rom";
defparam ram_block1a142.port_a_address_clear = "none";
defparam ram_block1a142.port_a_address_width = 13;
defparam ram_block1a142.port_a_data_out_clear = "none";
defparam ram_block1a142.port_a_data_out_clock = "clock0";
defparam ram_block1a142.port_a_data_width = 1;
defparam ram_block1a142.port_a_first_address = 40960;
defparam ram_block1a142.port_a_first_bit_number = 22;
defparam ram_block1a142.port_a_last_address = 49151;
defparam ram_block1a142.port_a_logical_ram_depth = 65536;
defparam ram_block1a142.port_a_logical_ram_width = 24;
defparam ram_block1a142.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a142.ram_block_type = "auto";
defparam ram_block1a142.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a142.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a142.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a142.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a166(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a166_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a166.clk0_core_clock_enable = "ena0";
defparam ram_block1a166.clk0_input_clock_enable = "ena0";
defparam ram_block1a166.clk0_output_clock_enable = "ena0";
defparam ram_block1a166.data_interleave_offset_in_bits = 1;
defparam ram_block1a166.data_interleave_width_in_bits = 1;
defparam ram_block1a166.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a166.init_file_layout = "port_a";
defparam ram_block1a166.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a166.operation_mode = "rom";
defparam ram_block1a166.port_a_address_clear = "none";
defparam ram_block1a166.port_a_address_width = 13;
defparam ram_block1a166.port_a_data_out_clear = "none";
defparam ram_block1a166.port_a_data_out_clock = "clock0";
defparam ram_block1a166.port_a_data_width = 1;
defparam ram_block1a166.port_a_first_address = 49152;
defparam ram_block1a166.port_a_first_bit_number = 22;
defparam ram_block1a166.port_a_last_address = 57343;
defparam ram_block1a166.port_a_logical_ram_depth = 65536;
defparam ram_block1a166.port_a_logical_ram_width = 24;
defparam ram_block1a166.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a166.ram_block_type = "auto";
defparam ram_block1a166.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a166.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a166.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a166.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a190(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a190_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a190.clk0_core_clock_enable = "ena0";
defparam ram_block1a190.clk0_input_clock_enable = "ena0";
defparam ram_block1a190.clk0_output_clock_enable = "ena0";
defparam ram_block1a190.data_interleave_offset_in_bits = 1;
defparam ram_block1a190.data_interleave_width_in_bits = 1;
defparam ram_block1a190.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a190.init_file_layout = "port_a";
defparam ram_block1a190.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a190.operation_mode = "rom";
defparam ram_block1a190.port_a_address_clear = "none";
defparam ram_block1a190.port_a_address_width = 13;
defparam ram_block1a190.port_a_data_out_clear = "none";
defparam ram_block1a190.port_a_data_out_clock = "clock0";
defparam ram_block1a190.port_a_data_width = 1;
defparam ram_block1a190.port_a_first_address = 57344;
defparam ram_block1a190.port_a_first_bit_number = 22;
defparam ram_block1a190.port_a_last_address = 65535;
defparam ram_block1a190.port_a_logical_ram_depth = 65536;
defparam ram_block1a190.port_a_logical_ram_width = 24;
defparam ram_block1a190.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a190.ram_block_type = "auto";
defparam ram_block1a190.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a190.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a190.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a190.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a70(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a70_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a70.clk0_core_clock_enable = "ena0";
defparam ram_block1a70.clk0_input_clock_enable = "ena0";
defparam ram_block1a70.clk0_output_clock_enable = "ena0";
defparam ram_block1a70.data_interleave_offset_in_bits = 1;
defparam ram_block1a70.data_interleave_width_in_bits = 1;
defparam ram_block1a70.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a70.init_file_layout = "port_a";
defparam ram_block1a70.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a70.operation_mode = "rom";
defparam ram_block1a70.port_a_address_clear = "none";
defparam ram_block1a70.port_a_address_width = 13;
defparam ram_block1a70.port_a_data_out_clear = "none";
defparam ram_block1a70.port_a_data_out_clock = "clock0";
defparam ram_block1a70.port_a_data_width = 1;
defparam ram_block1a70.port_a_first_address = 16384;
defparam ram_block1a70.port_a_first_bit_number = 22;
defparam ram_block1a70.port_a_last_address = 24575;
defparam ram_block1a70.port_a_logical_ram_depth = 65536;
defparam ram_block1a70.port_a_logical_ram_width = 24;
defparam ram_block1a70.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a70.ram_block_type = "auto";
defparam ram_block1a70.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a70.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a70.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a70.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a94(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a94_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a94.clk0_core_clock_enable = "ena0";
defparam ram_block1a94.clk0_input_clock_enable = "ena0";
defparam ram_block1a94.clk0_output_clock_enable = "ena0";
defparam ram_block1a94.data_interleave_offset_in_bits = 1;
defparam ram_block1a94.data_interleave_width_in_bits = 1;
defparam ram_block1a94.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a94.init_file_layout = "port_a";
defparam ram_block1a94.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a94.operation_mode = "rom";
defparam ram_block1a94.port_a_address_clear = "none";
defparam ram_block1a94.port_a_address_width = 13;
defparam ram_block1a94.port_a_data_out_clear = "none";
defparam ram_block1a94.port_a_data_out_clock = "clock0";
defparam ram_block1a94.port_a_data_width = 1;
defparam ram_block1a94.port_a_first_address = 24576;
defparam ram_block1a94.port_a_first_bit_number = 22;
defparam ram_block1a94.port_a_last_address = 32767;
defparam ram_block1a94.port_a_logical_ram_depth = 65536;
defparam ram_block1a94.port_a_logical_ram_width = 24;
defparam ram_block1a94.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a94.ram_block_type = "auto";
defparam ram_block1a94.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a94.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a94.mem_init1 = "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a94.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a22(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.clk0_output_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "rom";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "clock0";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 8191;
defparam ram_block1a22.port_a_logical_ram_depth = 65536;
defparam ram_block1a22.port_a_logical_ram_width = 24;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a22.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a46(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a46_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a46.clk0_core_clock_enable = "ena0";
defparam ram_block1a46.clk0_input_clock_enable = "ena0";
defparam ram_block1a46.clk0_output_clock_enable = "ena0";
defparam ram_block1a46.data_interleave_offset_in_bits = 1;
defparam ram_block1a46.data_interleave_width_in_bits = 1;
defparam ram_block1a46.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a46.init_file_layout = "port_a";
defparam ram_block1a46.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a46.operation_mode = "rom";
defparam ram_block1a46.port_a_address_clear = "none";
defparam ram_block1a46.port_a_address_width = 13;
defparam ram_block1a46.port_a_data_out_clear = "none";
defparam ram_block1a46.port_a_data_out_clock = "clock0";
defparam ram_block1a46.port_a_data_width = 1;
defparam ram_block1a46.port_a_first_address = 8192;
defparam ram_block1a46.port_a_first_bit_number = 22;
defparam ram_block1a46.port_a_last_address = 16383;
defparam ram_block1a46.port_a_logical_ram_depth = 65536;
defparam ram_block1a46.port_a_logical_ram_width = 24;
defparam ram_block1a46.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a46.ram_block_type = "auto";
defparam ram_block1a46.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a46.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a46.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a46.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a119(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a119_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a119.clk0_core_clock_enable = "ena0";
defparam ram_block1a119.clk0_input_clock_enable = "ena0";
defparam ram_block1a119.clk0_output_clock_enable = "ena0";
defparam ram_block1a119.data_interleave_offset_in_bits = 1;
defparam ram_block1a119.data_interleave_width_in_bits = 1;
defparam ram_block1a119.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a119.init_file_layout = "port_a";
defparam ram_block1a119.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a119.operation_mode = "rom";
defparam ram_block1a119.port_a_address_clear = "none";
defparam ram_block1a119.port_a_address_width = 13;
defparam ram_block1a119.port_a_data_out_clear = "none";
defparam ram_block1a119.port_a_data_out_clock = "clock0";
defparam ram_block1a119.port_a_data_width = 1;
defparam ram_block1a119.port_a_first_address = 32768;
defparam ram_block1a119.port_a_first_bit_number = 23;
defparam ram_block1a119.port_a_last_address = 40959;
defparam ram_block1a119.port_a_logical_ram_depth = 65536;
defparam ram_block1a119.port_a_logical_ram_width = 24;
defparam ram_block1a119.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a119.ram_block_type = "auto";
defparam ram_block1a119.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a119.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a119.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a119.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE";

cyclonev_ram_block ram_block1a143(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a143_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a143.clk0_core_clock_enable = "ena0";
defparam ram_block1a143.clk0_input_clock_enable = "ena0";
defparam ram_block1a143.clk0_output_clock_enable = "ena0";
defparam ram_block1a143.data_interleave_offset_in_bits = 1;
defparam ram_block1a143.data_interleave_width_in_bits = 1;
defparam ram_block1a143.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a143.init_file_layout = "port_a";
defparam ram_block1a143.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a143.operation_mode = "rom";
defparam ram_block1a143.port_a_address_clear = "none";
defparam ram_block1a143.port_a_address_width = 13;
defparam ram_block1a143.port_a_data_out_clear = "none";
defparam ram_block1a143.port_a_data_out_clock = "clock0";
defparam ram_block1a143.port_a_data_width = 1;
defparam ram_block1a143.port_a_first_address = 40960;
defparam ram_block1a143.port_a_first_bit_number = 23;
defparam ram_block1a143.port_a_last_address = 49151;
defparam ram_block1a143.port_a_logical_ram_depth = 65536;
defparam ram_block1a143.port_a_logical_ram_width = 24;
defparam ram_block1a143.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a143.ram_block_type = "auto";
defparam ram_block1a143.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a143.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a143.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a143.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a167(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a167_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a167.clk0_core_clock_enable = "ena0";
defparam ram_block1a167.clk0_input_clock_enable = "ena0";
defparam ram_block1a167.clk0_output_clock_enable = "ena0";
defparam ram_block1a167.data_interleave_offset_in_bits = 1;
defparam ram_block1a167.data_interleave_width_in_bits = 1;
defparam ram_block1a167.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a167.init_file_layout = "port_a";
defparam ram_block1a167.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a167.operation_mode = "rom";
defparam ram_block1a167.port_a_address_clear = "none";
defparam ram_block1a167.port_a_address_width = 13;
defparam ram_block1a167.port_a_data_out_clear = "none";
defparam ram_block1a167.port_a_data_out_clock = "clock0";
defparam ram_block1a167.port_a_data_width = 1;
defparam ram_block1a167.port_a_first_address = 49152;
defparam ram_block1a167.port_a_first_bit_number = 23;
defparam ram_block1a167.port_a_last_address = 57343;
defparam ram_block1a167.port_a_logical_ram_depth = 65536;
defparam ram_block1a167.port_a_logical_ram_width = 24;
defparam ram_block1a167.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a167.ram_block_type = "auto";
defparam ram_block1a167.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a167.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a167.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a167.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a191(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a191_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a191.clk0_core_clock_enable = "ena0";
defparam ram_block1a191.clk0_input_clock_enable = "ena0";
defparam ram_block1a191.clk0_output_clock_enable = "ena0";
defparam ram_block1a191.data_interleave_offset_in_bits = 1;
defparam ram_block1a191.data_interleave_width_in_bits = 1;
defparam ram_block1a191.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a191.init_file_layout = "port_a";
defparam ram_block1a191.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a191.operation_mode = "rom";
defparam ram_block1a191.port_a_address_clear = "none";
defparam ram_block1a191.port_a_address_width = 13;
defparam ram_block1a191.port_a_data_out_clear = "none";
defparam ram_block1a191.port_a_data_out_clock = "clock0";
defparam ram_block1a191.port_a_data_width = 1;
defparam ram_block1a191.port_a_first_address = 57344;
defparam ram_block1a191.port_a_first_bit_number = 23;
defparam ram_block1a191.port_a_last_address = 65535;
defparam ram_block1a191.port_a_logical_ram_depth = 65536;
defparam ram_block1a191.port_a_logical_ram_width = 24;
defparam ram_block1a191.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a191.ram_block_type = "auto";
defparam ram_block1a191.mem_init3 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a191.mem_init2 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a191.mem_init1 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
defparam ram_block1a191.mem_init0 = "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

cyclonev_ram_block ram_block1a71(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a71_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a71.clk0_core_clock_enable = "ena0";
defparam ram_block1a71.clk0_input_clock_enable = "ena0";
defparam ram_block1a71.clk0_output_clock_enable = "ena0";
defparam ram_block1a71.data_interleave_offset_in_bits = 1;
defparam ram_block1a71.data_interleave_width_in_bits = 1;
defparam ram_block1a71.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a71.init_file_layout = "port_a";
defparam ram_block1a71.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a71.operation_mode = "rom";
defparam ram_block1a71.port_a_address_clear = "none";
defparam ram_block1a71.port_a_address_width = 13;
defparam ram_block1a71.port_a_data_out_clear = "none";
defparam ram_block1a71.port_a_data_out_clock = "clock0";
defparam ram_block1a71.port_a_data_width = 1;
defparam ram_block1a71.port_a_first_address = 16384;
defparam ram_block1a71.port_a_first_bit_number = 23;
defparam ram_block1a71.port_a_last_address = 24575;
defparam ram_block1a71.port_a_logical_ram_depth = 65536;
defparam ram_block1a71.port_a_logical_ram_width = 24;
defparam ram_block1a71.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a71.ram_block_type = "auto";
defparam ram_block1a71.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a71.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a71.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a71.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a95(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a95_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a95.clk0_core_clock_enable = "ena0";
defparam ram_block1a95.clk0_input_clock_enable = "ena0";
defparam ram_block1a95.clk0_output_clock_enable = "ena0";
defparam ram_block1a95.data_interleave_offset_in_bits = 1;
defparam ram_block1a95.data_interleave_width_in_bits = 1;
defparam ram_block1a95.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a95.init_file_layout = "port_a";
defparam ram_block1a95.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a95.operation_mode = "rom";
defparam ram_block1a95.port_a_address_clear = "none";
defparam ram_block1a95.port_a_address_width = 13;
defparam ram_block1a95.port_a_data_out_clear = "none";
defparam ram_block1a95.port_a_data_out_clock = "clock0";
defparam ram_block1a95.port_a_data_width = 1;
defparam ram_block1a95.port_a_first_address = 24576;
defparam ram_block1a95.port_a_first_bit_number = 23;
defparam ram_block1a95.port_a_last_address = 32767;
defparam ram_block1a95.port_a_logical_ram_depth = 65536;
defparam ram_block1a95.port_a_logical_ram_width = 24;
defparam ram_block1a95.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a95.ram_block_type = "auto";
defparam ram_block1a95.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a95.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a95.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a95.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a23(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.clk0_output_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "rom";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "clock0";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 8191;
defparam ram_block1a23.port_a_logical_ram_depth = 65536;
defparam ram_block1a23.port_a_logical_ram_width = 24;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a47(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a47_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a47.clk0_core_clock_enable = "ena0";
defparam ram_block1a47.clk0_input_clock_enable = "ena0";
defparam ram_block1a47.clk0_output_clock_enable = "ena0";
defparam ram_block1a47.data_interleave_offset_in_bits = 1;
defparam ram_block1a47.data_interleave_width_in_bits = 1;
defparam ram_block1a47.init_file = "sine_nco_ii_0_sin.hex";
defparam ram_block1a47.init_file_layout = "port_a";
defparam ram_block1a47.logical_ram_name = "sine_nco_ii_0:nco_ii_0|asj_nco_as_m_cen:ux0120|altsyncram:altsyncram_component0|altsyncram_jtf1:auto_generated|ALTSYNCRAM";
defparam ram_block1a47.operation_mode = "rom";
defparam ram_block1a47.port_a_address_clear = "none";
defparam ram_block1a47.port_a_address_width = 13;
defparam ram_block1a47.port_a_data_out_clear = "none";
defparam ram_block1a47.port_a_data_out_clock = "clock0";
defparam ram_block1a47.port_a_data_width = 1;
defparam ram_block1a47.port_a_first_address = 8192;
defparam ram_block1a47.port_a_first_bit_number = 23;
defparam ram_block1a47.port_a_last_address = 16383;
defparam ram_block1a47.port_a_logical_ram_depth = 65536;
defparam ram_block1a47.port_a_logical_ram_width = 24;
defparam ram_block1a47.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a47.ram_block_type = "auto";
defparam ram_block1a47.mem_init3 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a47.mem_init2 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a47.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a47.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

dffeas \out_address_reg_a[2] (
	.clk(clock0),
	.d(\address_reg_a[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken0),
	.q(out_address_reg_a_2),
	.prn(vcc));
defparam \out_address_reg_a[2] .is_wysiwyg = "true";
defparam \out_address_reg_a[2] .power_up = "low";

dffeas \out_address_reg_a[0] (
	.clk(clock0),
	.d(\address_reg_a[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken0),
	.q(out_address_reg_a_0),
	.prn(vcc));
defparam \out_address_reg_a[0] .is_wysiwyg = "true";
defparam \out_address_reg_a[0] .power_up = "low";

dffeas \out_address_reg_a[1] (
	.clk(clock0),
	.d(\address_reg_a[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken0),
	.q(out_address_reg_a_1),
	.prn(vcc));
defparam \out_address_reg_a[1] .is_wysiwyg = "true";
defparam \out_address_reg_a[1] .power_up = "low";

dffeas \address_reg_a[2] (
	.clk(clock0),
	.d(address_a[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken0),
	.q(\address_reg_a[2]~q ),
	.prn(vcc));
defparam \address_reg_a[2] .is_wysiwyg = "true";
defparam \address_reg_a[2] .power_up = "low";

dffeas \address_reg_a[0] (
	.clk(clock0),
	.d(address_a[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken0),
	.q(\address_reg_a[0]~q ),
	.prn(vcc));
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";

dffeas \address_reg_a[1] (
	.clk(clock0),
	.d(address_a[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken0),
	.q(\address_reg_a[1]~q ),
	.prn(vcc));
defparam \address_reg_a[1] .is_wysiwyg = "true";
defparam \address_reg_a[1] .power_up = "low";

endmodule

module sine_asj_nco_fxx (
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_31,
	pipeline_dffe_15,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	clk,
	reset_n,
	clken,
	freq_mod_i_16,
	phi_inc_i_16,
	freq_mod_i_17,
	phi_inc_i_17,
	freq_mod_i_18,
	phi_inc_i_18,
	freq_mod_i_19,
	phi_inc_i_19,
	freq_mod_i_20,
	phi_inc_i_20,
	freq_mod_i_21,
	phi_inc_i_21,
	freq_mod_i_22,
	phi_inc_i_22,
	freq_mod_i_23,
	phi_inc_i_23,
	freq_mod_i_24,
	phi_inc_i_24,
	freq_mod_i_25,
	phi_inc_i_25,
	freq_mod_i_26,
	phi_inc_i_26,
	freq_mod_i_27,
	phi_inc_i_27,
	freq_mod_i_28,
	phi_inc_i_28,
	freq_mod_i_31,
	phi_inc_i_31,
	freq_mod_i_15,
	phi_inc_i_15,
	freq_mod_i_29,
	phi_inc_i_29,
	freq_mod_i_30,
	phi_inc_i_30,
	freq_mod_i_14,
	phi_inc_i_14,
	freq_mod_i_13,
	phi_inc_i_13,
	freq_mod_i_12,
	phi_inc_i_12,
	freq_mod_i_11,
	phi_inc_i_11,
	freq_mod_i_10,
	phi_inc_i_10,
	freq_mod_i_9,
	phi_inc_i_9,
	freq_mod_i_8,
	phi_inc_i_8,
	freq_mod_i_7,
	phi_inc_i_7,
	freq_mod_i_6,
	phi_inc_i_6,
	freq_mod_i_5,
	phi_inc_i_5,
	freq_mod_i_4,
	phi_inc_i_4,
	freq_mod_i_3,
	phi_inc_i_3,
	freq_mod_i_2,
	phi_inc_i_2,
	freq_mod_i_1,
	phi_inc_i_1,
	freq_mod_i_0,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_31;
output 	pipeline_dffe_15;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
input 	clk;
input 	reset_n;
input 	clken;
input 	freq_mod_i_16;
input 	phi_inc_i_16;
input 	freq_mod_i_17;
input 	phi_inc_i_17;
input 	freq_mod_i_18;
input 	phi_inc_i_18;
input 	freq_mod_i_19;
input 	phi_inc_i_19;
input 	freq_mod_i_20;
input 	phi_inc_i_20;
input 	freq_mod_i_21;
input 	phi_inc_i_21;
input 	freq_mod_i_22;
input 	phi_inc_i_22;
input 	freq_mod_i_23;
input 	phi_inc_i_23;
input 	freq_mod_i_24;
input 	phi_inc_i_24;
input 	freq_mod_i_25;
input 	phi_inc_i_25;
input 	freq_mod_i_26;
input 	phi_inc_i_26;
input 	freq_mod_i_27;
input 	phi_inc_i_27;
input 	freq_mod_i_28;
input 	phi_inc_i_28;
input 	freq_mod_i_31;
input 	phi_inc_i_31;
input 	freq_mod_i_15;
input 	phi_inc_i_15;
input 	freq_mod_i_29;
input 	phi_inc_i_29;
input 	freq_mod_i_30;
input 	phi_inc_i_30;
input 	freq_mod_i_14;
input 	phi_inc_i_14;
input 	freq_mod_i_13;
input 	phi_inc_i_13;
input 	freq_mod_i_12;
input 	phi_inc_i_12;
input 	freq_mod_i_11;
input 	phi_inc_i_11;
input 	freq_mod_i_10;
input 	phi_inc_i_10;
input 	freq_mod_i_9;
input 	phi_inc_i_9;
input 	freq_mod_i_8;
input 	phi_inc_i_8;
input 	freq_mod_i_7;
input 	phi_inc_i_7;
input 	freq_mod_i_6;
input 	phi_inc_i_6;
input 	freq_mod_i_5;
input 	phi_inc_i_5;
input 	freq_mod_i_4;
input 	phi_inc_i_4;
input 	freq_mod_i_3;
input 	phi_inc_i_3;
input 	freq_mod_i_2;
input 	phi_inc_i_2;
input 	freq_mod_i_1;
input 	phi_inc_i_1;
input 	freq_mod_i_0;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_lpm_add_sub_2 acc(
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken),
	.freq_mod_i_16(freq_mod_i_16),
	.phi_inc_i_16(phi_inc_i_16),
	.freq_mod_i_17(freq_mod_i_17),
	.phi_inc_i_17(phi_inc_i_17),
	.freq_mod_i_18(freq_mod_i_18),
	.phi_inc_i_18(phi_inc_i_18),
	.freq_mod_i_19(freq_mod_i_19),
	.phi_inc_i_19(phi_inc_i_19),
	.freq_mod_i_20(freq_mod_i_20),
	.phi_inc_i_20(phi_inc_i_20),
	.freq_mod_i_21(freq_mod_i_21),
	.phi_inc_i_21(phi_inc_i_21),
	.freq_mod_i_22(freq_mod_i_22),
	.phi_inc_i_22(phi_inc_i_22),
	.freq_mod_i_23(freq_mod_i_23),
	.phi_inc_i_23(phi_inc_i_23),
	.freq_mod_i_24(freq_mod_i_24),
	.phi_inc_i_24(phi_inc_i_24),
	.freq_mod_i_25(freq_mod_i_25),
	.phi_inc_i_25(phi_inc_i_25),
	.freq_mod_i_26(freq_mod_i_26),
	.phi_inc_i_26(phi_inc_i_26),
	.freq_mod_i_27(freq_mod_i_27),
	.phi_inc_i_27(phi_inc_i_27),
	.freq_mod_i_28(freq_mod_i_28),
	.phi_inc_i_28(phi_inc_i_28),
	.freq_mod_i_31(freq_mod_i_31),
	.phi_inc_i_31(phi_inc_i_31),
	.freq_mod_i_15(freq_mod_i_15),
	.phi_inc_i_15(phi_inc_i_15),
	.freq_mod_i_29(freq_mod_i_29),
	.phi_inc_i_29(phi_inc_i_29),
	.freq_mod_i_30(freq_mod_i_30),
	.phi_inc_i_30(phi_inc_i_30),
	.freq_mod_i_14(freq_mod_i_14),
	.phi_inc_i_14(phi_inc_i_14),
	.freq_mod_i_13(freq_mod_i_13),
	.phi_inc_i_13(phi_inc_i_13),
	.freq_mod_i_12(freq_mod_i_12),
	.phi_inc_i_12(phi_inc_i_12),
	.freq_mod_i_11(freq_mod_i_11),
	.phi_inc_i_11(phi_inc_i_11),
	.freq_mod_i_10(freq_mod_i_10),
	.phi_inc_i_10(phi_inc_i_10),
	.freq_mod_i_9(freq_mod_i_9),
	.phi_inc_i_9(phi_inc_i_9),
	.freq_mod_i_8(freq_mod_i_8),
	.phi_inc_i_8(phi_inc_i_8),
	.freq_mod_i_7(freq_mod_i_7),
	.phi_inc_i_7(phi_inc_i_7),
	.freq_mod_i_6(freq_mod_i_6),
	.phi_inc_i_6(phi_inc_i_6),
	.freq_mod_i_5(freq_mod_i_5),
	.phi_inc_i_5(phi_inc_i_5),
	.freq_mod_i_4(freq_mod_i_4),
	.phi_inc_i_4(phi_inc_i_4),
	.freq_mod_i_3(freq_mod_i_3),
	.phi_inc_i_3(phi_inc_i_3),
	.freq_mod_i_2(freq_mod_i_2),
	.phi_inc_i_2(phi_inc_i_2),
	.freq_mod_i_1(freq_mod_i_1),
	.phi_inc_i_1(phi_inc_i_1),
	.freq_mod_i_0(freq_mod_i_0),
	.phi_inc_i_0(phi_inc_i_0));

endmodule

module sine_lpm_add_sub_2 (
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_31,
	pipeline_dffe_15,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	clock,
	reset_n,
	clken,
	freq_mod_i_16,
	phi_inc_i_16,
	freq_mod_i_17,
	phi_inc_i_17,
	freq_mod_i_18,
	phi_inc_i_18,
	freq_mod_i_19,
	phi_inc_i_19,
	freq_mod_i_20,
	phi_inc_i_20,
	freq_mod_i_21,
	phi_inc_i_21,
	freq_mod_i_22,
	phi_inc_i_22,
	freq_mod_i_23,
	phi_inc_i_23,
	freq_mod_i_24,
	phi_inc_i_24,
	freq_mod_i_25,
	phi_inc_i_25,
	freq_mod_i_26,
	phi_inc_i_26,
	freq_mod_i_27,
	phi_inc_i_27,
	freq_mod_i_28,
	phi_inc_i_28,
	freq_mod_i_31,
	phi_inc_i_31,
	freq_mod_i_15,
	phi_inc_i_15,
	freq_mod_i_29,
	phi_inc_i_29,
	freq_mod_i_30,
	phi_inc_i_30,
	freq_mod_i_14,
	phi_inc_i_14,
	freq_mod_i_13,
	phi_inc_i_13,
	freq_mod_i_12,
	phi_inc_i_12,
	freq_mod_i_11,
	phi_inc_i_11,
	freq_mod_i_10,
	phi_inc_i_10,
	freq_mod_i_9,
	phi_inc_i_9,
	freq_mod_i_8,
	phi_inc_i_8,
	freq_mod_i_7,
	phi_inc_i_7,
	freq_mod_i_6,
	phi_inc_i_6,
	freq_mod_i_5,
	phi_inc_i_5,
	freq_mod_i_4,
	phi_inc_i_4,
	freq_mod_i_3,
	phi_inc_i_3,
	freq_mod_i_2,
	phi_inc_i_2,
	freq_mod_i_1,
	phi_inc_i_1,
	freq_mod_i_0,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_31;
output 	pipeline_dffe_15;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
input 	clock;
input 	reset_n;
input 	clken;
input 	freq_mod_i_16;
input 	phi_inc_i_16;
input 	freq_mod_i_17;
input 	phi_inc_i_17;
input 	freq_mod_i_18;
input 	phi_inc_i_18;
input 	freq_mod_i_19;
input 	phi_inc_i_19;
input 	freq_mod_i_20;
input 	phi_inc_i_20;
input 	freq_mod_i_21;
input 	phi_inc_i_21;
input 	freq_mod_i_22;
input 	phi_inc_i_22;
input 	freq_mod_i_23;
input 	phi_inc_i_23;
input 	freq_mod_i_24;
input 	phi_inc_i_24;
input 	freq_mod_i_25;
input 	phi_inc_i_25;
input 	freq_mod_i_26;
input 	phi_inc_i_26;
input 	freq_mod_i_27;
input 	phi_inc_i_27;
input 	freq_mod_i_28;
input 	phi_inc_i_28;
input 	freq_mod_i_31;
input 	phi_inc_i_31;
input 	freq_mod_i_15;
input 	phi_inc_i_15;
input 	freq_mod_i_29;
input 	phi_inc_i_29;
input 	freq_mod_i_30;
input 	phi_inc_i_30;
input 	freq_mod_i_14;
input 	phi_inc_i_14;
input 	freq_mod_i_13;
input 	phi_inc_i_13;
input 	freq_mod_i_12;
input 	phi_inc_i_12;
input 	freq_mod_i_11;
input 	phi_inc_i_11;
input 	freq_mod_i_10;
input 	phi_inc_i_10;
input 	freq_mod_i_9;
input 	phi_inc_i_9;
input 	freq_mod_i_8;
input 	phi_inc_i_8;
input 	freq_mod_i_7;
input 	phi_inc_i_7;
input 	freq_mod_i_6;
input 	phi_inc_i_6;
input 	freq_mod_i_5;
input 	phi_inc_i_5;
input 	freq_mod_i_4;
input 	phi_inc_i_4;
input 	freq_mod_i_3;
input 	phi_inc_i_3;
input 	freq_mod_i_2;
input 	phi_inc_i_2;
input 	freq_mod_i_1;
input 	phi_inc_i_1;
input 	freq_mod_i_0;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_add_sub_q0h auto_generated(
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken),
	.freq_mod_i_16(freq_mod_i_16),
	.phi_inc_i_16(phi_inc_i_16),
	.freq_mod_i_17(freq_mod_i_17),
	.phi_inc_i_17(phi_inc_i_17),
	.freq_mod_i_18(freq_mod_i_18),
	.phi_inc_i_18(phi_inc_i_18),
	.freq_mod_i_19(freq_mod_i_19),
	.phi_inc_i_19(phi_inc_i_19),
	.freq_mod_i_20(freq_mod_i_20),
	.phi_inc_i_20(phi_inc_i_20),
	.freq_mod_i_21(freq_mod_i_21),
	.phi_inc_i_21(phi_inc_i_21),
	.freq_mod_i_22(freq_mod_i_22),
	.phi_inc_i_22(phi_inc_i_22),
	.freq_mod_i_23(freq_mod_i_23),
	.phi_inc_i_23(phi_inc_i_23),
	.freq_mod_i_24(freq_mod_i_24),
	.phi_inc_i_24(phi_inc_i_24),
	.freq_mod_i_25(freq_mod_i_25),
	.phi_inc_i_25(phi_inc_i_25),
	.freq_mod_i_26(freq_mod_i_26),
	.phi_inc_i_26(phi_inc_i_26),
	.freq_mod_i_27(freq_mod_i_27),
	.phi_inc_i_27(phi_inc_i_27),
	.freq_mod_i_28(freq_mod_i_28),
	.phi_inc_i_28(phi_inc_i_28),
	.freq_mod_i_31(freq_mod_i_31),
	.phi_inc_i_31(phi_inc_i_31),
	.freq_mod_i_15(freq_mod_i_15),
	.phi_inc_i_15(phi_inc_i_15),
	.freq_mod_i_29(freq_mod_i_29),
	.phi_inc_i_29(phi_inc_i_29),
	.freq_mod_i_30(freq_mod_i_30),
	.phi_inc_i_30(phi_inc_i_30),
	.freq_mod_i_14(freq_mod_i_14),
	.phi_inc_i_14(phi_inc_i_14),
	.freq_mod_i_13(freq_mod_i_13),
	.phi_inc_i_13(phi_inc_i_13),
	.freq_mod_i_12(freq_mod_i_12),
	.phi_inc_i_12(phi_inc_i_12),
	.freq_mod_i_11(freq_mod_i_11),
	.phi_inc_i_11(phi_inc_i_11),
	.freq_mod_i_10(freq_mod_i_10),
	.phi_inc_i_10(phi_inc_i_10),
	.freq_mod_i_9(freq_mod_i_9),
	.phi_inc_i_9(phi_inc_i_9),
	.freq_mod_i_8(freq_mod_i_8),
	.phi_inc_i_8(phi_inc_i_8),
	.freq_mod_i_7(freq_mod_i_7),
	.phi_inc_i_7(phi_inc_i_7),
	.freq_mod_i_6(freq_mod_i_6),
	.phi_inc_i_6(phi_inc_i_6),
	.freq_mod_i_5(freq_mod_i_5),
	.phi_inc_i_5(phi_inc_i_5),
	.freq_mod_i_4(freq_mod_i_4),
	.phi_inc_i_4(phi_inc_i_4),
	.freq_mod_i_3(freq_mod_i_3),
	.phi_inc_i_3(phi_inc_i_3),
	.freq_mod_i_2(freq_mod_i_2),
	.phi_inc_i_2(phi_inc_i_2),
	.freq_mod_i_1(freq_mod_i_1),
	.phi_inc_i_1(phi_inc_i_1),
	.freq_mod_i_0(freq_mod_i_0),
	.phi_inc_i_0(phi_inc_i_0));

endmodule

module sine_add_sub_q0h (
	pipeline_dffe_16,
	pipeline_dffe_17,
	pipeline_dffe_18,
	pipeline_dffe_19,
	pipeline_dffe_20,
	pipeline_dffe_21,
	pipeline_dffe_22,
	pipeline_dffe_23,
	pipeline_dffe_24,
	pipeline_dffe_25,
	pipeline_dffe_26,
	pipeline_dffe_27,
	pipeline_dffe_28,
	pipeline_dffe_31,
	pipeline_dffe_15,
	pipeline_dffe_29,
	pipeline_dffe_30,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	clock,
	reset_n,
	clken,
	freq_mod_i_16,
	phi_inc_i_16,
	freq_mod_i_17,
	phi_inc_i_17,
	freq_mod_i_18,
	phi_inc_i_18,
	freq_mod_i_19,
	phi_inc_i_19,
	freq_mod_i_20,
	phi_inc_i_20,
	freq_mod_i_21,
	phi_inc_i_21,
	freq_mod_i_22,
	phi_inc_i_22,
	freq_mod_i_23,
	phi_inc_i_23,
	freq_mod_i_24,
	phi_inc_i_24,
	freq_mod_i_25,
	phi_inc_i_25,
	freq_mod_i_26,
	phi_inc_i_26,
	freq_mod_i_27,
	phi_inc_i_27,
	freq_mod_i_28,
	phi_inc_i_28,
	freq_mod_i_31,
	phi_inc_i_31,
	freq_mod_i_15,
	phi_inc_i_15,
	freq_mod_i_29,
	phi_inc_i_29,
	freq_mod_i_30,
	phi_inc_i_30,
	freq_mod_i_14,
	phi_inc_i_14,
	freq_mod_i_13,
	phi_inc_i_13,
	freq_mod_i_12,
	phi_inc_i_12,
	freq_mod_i_11,
	phi_inc_i_11,
	freq_mod_i_10,
	phi_inc_i_10,
	freq_mod_i_9,
	phi_inc_i_9,
	freq_mod_i_8,
	phi_inc_i_8,
	freq_mod_i_7,
	phi_inc_i_7,
	freq_mod_i_6,
	phi_inc_i_6,
	freq_mod_i_5,
	phi_inc_i_5,
	freq_mod_i_4,
	phi_inc_i_4,
	freq_mod_i_3,
	phi_inc_i_3,
	freq_mod_i_2,
	phi_inc_i_2,
	freq_mod_i_1,
	phi_inc_i_1,
	freq_mod_i_0,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
output 	pipeline_dffe_18;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
output 	pipeline_dffe_21;
output 	pipeline_dffe_22;
output 	pipeline_dffe_23;
output 	pipeline_dffe_24;
output 	pipeline_dffe_25;
output 	pipeline_dffe_26;
output 	pipeline_dffe_27;
output 	pipeline_dffe_28;
output 	pipeline_dffe_31;
output 	pipeline_dffe_15;
output 	pipeline_dffe_29;
output 	pipeline_dffe_30;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
input 	clock;
input 	reset_n;
input 	clken;
input 	freq_mod_i_16;
input 	phi_inc_i_16;
input 	freq_mod_i_17;
input 	phi_inc_i_17;
input 	freq_mod_i_18;
input 	phi_inc_i_18;
input 	freq_mod_i_19;
input 	phi_inc_i_19;
input 	freq_mod_i_20;
input 	phi_inc_i_20;
input 	freq_mod_i_21;
input 	phi_inc_i_21;
input 	freq_mod_i_22;
input 	phi_inc_i_22;
input 	freq_mod_i_23;
input 	phi_inc_i_23;
input 	freq_mod_i_24;
input 	phi_inc_i_24;
input 	freq_mod_i_25;
input 	phi_inc_i_25;
input 	freq_mod_i_26;
input 	phi_inc_i_26;
input 	freq_mod_i_27;
input 	phi_inc_i_27;
input 	freq_mod_i_28;
input 	phi_inc_i_28;
input 	freq_mod_i_31;
input 	phi_inc_i_31;
input 	freq_mod_i_15;
input 	phi_inc_i_15;
input 	freq_mod_i_29;
input 	phi_inc_i_29;
input 	freq_mod_i_30;
input 	phi_inc_i_30;
input 	freq_mod_i_14;
input 	phi_inc_i_14;
input 	freq_mod_i_13;
input 	phi_inc_i_13;
input 	freq_mod_i_12;
input 	phi_inc_i_12;
input 	freq_mod_i_11;
input 	phi_inc_i_11;
input 	freq_mod_i_10;
input 	phi_inc_i_10;
input 	freq_mod_i_9;
input 	phi_inc_i_9;
input 	freq_mod_i_8;
input 	phi_inc_i_8;
input 	freq_mod_i_7;
input 	phi_inc_i_7;
input 	freq_mod_i_6;
input 	phi_inc_i_6;
input 	freq_mod_i_5;
input 	phi_inc_i_5;
input 	freq_mod_i_4;
input 	phi_inc_i_4;
input 	freq_mod_i_3;
input 	phi_inc_i_3;
input 	freq_mod_i_2;
input 	phi_inc_i_2;
input 	freq_mod_i_1;
input 	phi_inc_i_1;
input 	freq_mod_i_0;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~126 ;
wire \op_1~122 ;
wire \op_1~118 ;
wire \op_1~114 ;
wire \op_1~110 ;
wire \op_1~106 ;
wire \op_1~102 ;
wire \op_1~98 ;
wire \op_1~94 ;
wire \op_1~90 ;
wire \op_1~86 ;
wire \op_1~82 ;
wire \op_1~78 ;
wire \op_1~74 ;
wire \op_1~70 ;
wire \op_1~58 ;
wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~6 ;
wire \op_1~9_sumout ;
wire \op_1~10 ;
wire \op_1~13_sumout ;
wire \op_1~14 ;
wire \op_1~17_sumout ;
wire \op_1~18 ;
wire \op_1~21_sumout ;
wire \op_1~22 ;
wire \op_1~25_sumout ;
wire \op_1~26 ;
wire \op_1~29_sumout ;
wire \op_1~30 ;
wire \op_1~33_sumout ;
wire \op_1~34 ;
wire \op_1~37_sumout ;
wire \op_1~38 ;
wire \op_1~41_sumout ;
wire \op_1~42 ;
wire \op_1~45_sumout ;
wire \op_1~46 ;
wire \op_1~49_sumout ;
wire \op_1~50 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~73_sumout ;
wire \op_1~77_sumout ;
wire \op_1~81_sumout ;
wire \op_1~85_sumout ;
wire \op_1~89_sumout ;
wire \op_1~93_sumout ;
wire \op_1~97_sumout ;
wire \op_1~101_sumout ;
wire \op_1~105_sumout ;
wire \op_1~109_sumout ;
wire \op_1~113_sumout ;
wire \op_1~117_sumout ;
wire \op_1~121_sumout ;
wire \op_1~125_sumout ;


dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[18] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \pipeline_dffe[18] .is_wysiwyg = "true";
defparam \pipeline_dffe[18] .power_up = "low";

dffeas \pipeline_dffe[19] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \pipeline_dffe[19] .is_wysiwyg = "true";
defparam \pipeline_dffe[19] .power_up = "low";

dffeas \pipeline_dffe[20] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_20),
	.prn(vcc));
defparam \pipeline_dffe[20] .is_wysiwyg = "true";
defparam \pipeline_dffe[20] .power_up = "low";

dffeas \pipeline_dffe[21] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_21),
	.prn(vcc));
defparam \pipeline_dffe[21] .is_wysiwyg = "true";
defparam \pipeline_dffe[21] .power_up = "low";

dffeas \pipeline_dffe[22] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_22),
	.prn(vcc));
defparam \pipeline_dffe[22] .is_wysiwyg = "true";
defparam \pipeline_dffe[22] .power_up = "low";

dffeas \pipeline_dffe[23] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_23),
	.prn(vcc));
defparam \pipeline_dffe[23] .is_wysiwyg = "true";
defparam \pipeline_dffe[23] .power_up = "low";

dffeas \pipeline_dffe[24] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_24),
	.prn(vcc));
defparam \pipeline_dffe[24] .is_wysiwyg = "true";
defparam \pipeline_dffe[24] .power_up = "low";

dffeas \pipeline_dffe[25] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_25),
	.prn(vcc));
defparam \pipeline_dffe[25] .is_wysiwyg = "true";
defparam \pipeline_dffe[25] .power_up = "low";

dffeas \pipeline_dffe[26] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_26),
	.prn(vcc));
defparam \pipeline_dffe[26] .is_wysiwyg = "true";
defparam \pipeline_dffe[26] .power_up = "low";

dffeas \pipeline_dffe[27] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_27),
	.prn(vcc));
defparam \pipeline_dffe[27] .is_wysiwyg = "true";
defparam \pipeline_dffe[27] .power_up = "low";

dffeas \pipeline_dffe[28] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_28),
	.prn(vcc));
defparam \pipeline_dffe[28] .is_wysiwyg = "true";
defparam \pipeline_dffe[28] .power_up = "low";

dffeas \pipeline_dffe[31] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_31),
	.prn(vcc));
defparam \pipeline_dffe[31] .is_wysiwyg = "true";
defparam \pipeline_dffe[31] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[29] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_29),
	.prn(vcc));
defparam \pipeline_dffe[29] .is_wysiwyg = "true";
defparam \pipeline_dffe[29] .power_up = "low";

dffeas \pipeline_dffe[30] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_30),
	.prn(vcc));
defparam \pipeline_dffe[30] .is_wysiwyg = "true";
defparam \pipeline_dffe[30] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~73_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~77_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~81_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~85_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~89_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~93_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~97_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~101_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~105_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~109_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~113_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~117_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~121_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~125_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

cyclonev_lcell_comb \op_1~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_0),
	.datae(gnd),
	.dataf(!phi_inc_i_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~125_sumout ),
	.cout(\op_1~126 ),
	.shareout());
defparam \op_1~125 .extended_lut = "off";
defparam \op_1~125 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~125 .shared_arith = "off";

cyclonev_lcell_comb \op_1~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_1),
	.datae(gnd),
	.dataf(!phi_inc_i_1),
	.datag(gnd),
	.cin(\op_1~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~121_sumout ),
	.cout(\op_1~122 ),
	.shareout());
defparam \op_1~121 .extended_lut = "off";
defparam \op_1~121 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~121 .shared_arith = "off";

cyclonev_lcell_comb \op_1~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_2),
	.datae(gnd),
	.dataf(!phi_inc_i_2),
	.datag(gnd),
	.cin(\op_1~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~117_sumout ),
	.cout(\op_1~118 ),
	.shareout());
defparam \op_1~117 .extended_lut = "off";
defparam \op_1~117 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~117 .shared_arith = "off";

cyclonev_lcell_comb \op_1~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_3),
	.datae(gnd),
	.dataf(!phi_inc_i_3),
	.datag(gnd),
	.cin(\op_1~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~113_sumout ),
	.cout(\op_1~114 ),
	.shareout());
defparam \op_1~113 .extended_lut = "off";
defparam \op_1~113 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~113 .shared_arith = "off";

cyclonev_lcell_comb \op_1~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_4),
	.datae(gnd),
	.dataf(!phi_inc_i_4),
	.datag(gnd),
	.cin(\op_1~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~109_sumout ),
	.cout(\op_1~110 ),
	.shareout());
defparam \op_1~109 .extended_lut = "off";
defparam \op_1~109 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~109 .shared_arith = "off";

cyclonev_lcell_comb \op_1~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_5),
	.datae(gnd),
	.dataf(!phi_inc_i_5),
	.datag(gnd),
	.cin(\op_1~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~105_sumout ),
	.cout(\op_1~106 ),
	.shareout());
defparam \op_1~105 .extended_lut = "off";
defparam \op_1~105 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~105 .shared_arith = "off";

cyclonev_lcell_comb \op_1~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_6),
	.datae(gnd),
	.dataf(!phi_inc_i_6),
	.datag(gnd),
	.cin(\op_1~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~101_sumout ),
	.cout(\op_1~102 ),
	.shareout());
defparam \op_1~101 .extended_lut = "off";
defparam \op_1~101 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~101 .shared_arith = "off";

cyclonev_lcell_comb \op_1~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_7),
	.datae(gnd),
	.dataf(!phi_inc_i_7),
	.datag(gnd),
	.cin(\op_1~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~97_sumout ),
	.cout(\op_1~98 ),
	.shareout());
defparam \op_1~97 .extended_lut = "off";
defparam \op_1~97 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~97 .shared_arith = "off";

cyclonev_lcell_comb \op_1~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_8),
	.datae(gnd),
	.dataf(!phi_inc_i_8),
	.datag(gnd),
	.cin(\op_1~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~93_sumout ),
	.cout(\op_1~94 ),
	.shareout());
defparam \op_1~93 .extended_lut = "off";
defparam \op_1~93 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~93 .shared_arith = "off";

cyclonev_lcell_comb \op_1~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_9),
	.datae(gnd),
	.dataf(!phi_inc_i_9),
	.datag(gnd),
	.cin(\op_1~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~89_sumout ),
	.cout(\op_1~90 ),
	.shareout());
defparam \op_1~89 .extended_lut = "off";
defparam \op_1~89 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~89 .shared_arith = "off";

cyclonev_lcell_comb \op_1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_10),
	.datae(gnd),
	.dataf(!phi_inc_i_10),
	.datag(gnd),
	.cin(\op_1~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~85_sumout ),
	.cout(\op_1~86 ),
	.shareout());
defparam \op_1~85 .extended_lut = "off";
defparam \op_1~85 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~85 .shared_arith = "off";

cyclonev_lcell_comb \op_1~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_11),
	.datae(gnd),
	.dataf(!phi_inc_i_11),
	.datag(gnd),
	.cin(\op_1~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~81_sumout ),
	.cout(\op_1~82 ),
	.shareout());
defparam \op_1~81 .extended_lut = "off";
defparam \op_1~81 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~81 .shared_arith = "off";

cyclonev_lcell_comb \op_1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_12),
	.datae(gnd),
	.dataf(!phi_inc_i_12),
	.datag(gnd),
	.cin(\op_1~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~77_sumout ),
	.cout(\op_1~78 ),
	.shareout());
defparam \op_1~77 .extended_lut = "off";
defparam \op_1~77 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~77 .shared_arith = "off";

cyclonev_lcell_comb \op_1~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_13),
	.datae(gnd),
	.dataf(!phi_inc_i_13),
	.datag(gnd),
	.cin(\op_1~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~73_sumout ),
	.cout(\op_1~74 ),
	.shareout());
defparam \op_1~73 .extended_lut = "off";
defparam \op_1~73 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~73 .shared_arith = "off";

cyclonev_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_14),
	.datae(gnd),
	.dataf(!phi_inc_i_14),
	.datag(gnd),
	.cin(\op_1~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

cyclonev_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_15),
	.datae(gnd),
	.dataf(!phi_inc_i_15),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_16),
	.datae(gnd),
	.dataf(!phi_inc_i_16),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_17),
	.datae(gnd),
	.dataf(!phi_inc_i_17),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_18),
	.datae(gnd),
	.dataf(!phi_inc_i_18),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_19),
	.datae(gnd),
	.dataf(!phi_inc_i_19),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_20),
	.datae(gnd),
	.dataf(!phi_inc_i_20),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_21),
	.datae(gnd),
	.dataf(!phi_inc_i_21),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_22),
	.datae(gnd),
	.dataf(!phi_inc_i_22),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_23),
	.datae(gnd),
	.dataf(!phi_inc_i_23),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_24),
	.datae(gnd),
	.dataf(!phi_inc_i_24),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_25),
	.datae(gnd),
	.dataf(!phi_inc_i_25),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_26),
	.datae(gnd),
	.dataf(!phi_inc_i_26),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_27),
	.datae(gnd),
	.dataf(!phi_inc_i_27),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_28),
	.datae(gnd),
	.dataf(!phi_inc_i_28),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

cyclonev_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_29),
	.datae(gnd),
	.dataf(!phi_inc_i_29),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

cyclonev_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_30),
	.datae(gnd),
	.dataf(!phi_inc_i_30),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

cyclonev_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!freq_mod_i_31),
	.datae(gnd),
	.dataf(!phi_inc_i_31),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

endmodule

module sine_asj_nco_isdr (
	data_ready1,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	data_ready1;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lpm_counter_component|auto_generated|counter_reg_bit[3]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[2]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[1]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[0]~q ;
wire \data_ready~0_combout ;


sine_lpm_counter_1 lpm_counter_component(
	.counter_reg_bit_3(\lpm_counter_component|auto_generated|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\lpm_counter_component|auto_generated|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\lpm_counter_component|auto_generated|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\lpm_counter_component|auto_generated|counter_reg_bit[0]~q ),
	.clock(clk),
	.sclr(reset_n),
	.clken(clken));

dffeas data_ready(
	.clk(clk),
	.d(\data_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(data_ready1),
	.prn(vcc));
defparam data_ready.is_wysiwyg = "true";
defparam data_ready.power_up = "low";

cyclonev_lcell_comb \data_ready~0 (
	.dataa(!data_ready1),
	.datab(!clken),
	.datac(!\lpm_counter_component|auto_generated|counter_reg_bit[3]~q ),
	.datad(!\lpm_counter_component|auto_generated|counter_reg_bit[2]~q ),
	.datae(!\lpm_counter_component|auto_generated|counter_reg_bit[1]~q ),
	.dataf(!\lpm_counter_component|auto_generated|counter_reg_bit[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_ready~0 .extended_lut = "off";
defparam \data_ready~0 .lut_mask = 64'hFFFFFFFFFFFFFF7F;
defparam \data_ready~0 .shared_arith = "off";

endmodule

module sine_lpm_counter_1 (
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	clock,
	sclr,
	clken)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	clock;
input 	sclr;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_cntr_ski auto_generated(
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.clock(clock),
	.sclr(sclr),
	.clken(clken));

endmodule

module sine_cntr_ski (
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	clock,
	sclr,
	clken)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	clock;
input 	sclr;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita0~sumout ;


dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

endmodule

module sine_asj_nco_mob_rw (
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	data_out_10,
	data_out_11,
	data_out_12,
	data_out_13,
	data_out_14,
	data_out_15,
	data_out_16,
	data_out_17,
	data_out_18,
	data_out_19,
	data_out_20,
	data_out_21,
	data_out_22,
	data_out_23,
	ram_block1a96,
	ram_block1a120,
	ram_block1a144,
	ram_block1a168,
	ram_block1a48,
	ram_block1a72,
	ram_block1a0,
	ram_block1a24,
	ram_block1a97,
	ram_block1a121,
	ram_block1a145,
	ram_block1a169,
	ram_block1a49,
	ram_block1a73,
	ram_block1a1,
	ram_block1a25,
	ram_block1a98,
	ram_block1a122,
	ram_block1a146,
	ram_block1a170,
	ram_block1a50,
	ram_block1a74,
	ram_block1a2,
	ram_block1a26,
	ram_block1a99,
	ram_block1a123,
	ram_block1a147,
	ram_block1a171,
	ram_block1a51,
	ram_block1a75,
	ram_block1a3,
	ram_block1a27,
	ram_block1a100,
	ram_block1a124,
	ram_block1a148,
	ram_block1a172,
	ram_block1a52,
	ram_block1a76,
	ram_block1a4,
	ram_block1a28,
	ram_block1a101,
	ram_block1a125,
	ram_block1a149,
	ram_block1a173,
	ram_block1a53,
	ram_block1a77,
	ram_block1a5,
	ram_block1a29,
	ram_block1a102,
	ram_block1a126,
	ram_block1a150,
	ram_block1a174,
	ram_block1a54,
	ram_block1a78,
	ram_block1a6,
	ram_block1a30,
	ram_block1a103,
	ram_block1a127,
	ram_block1a151,
	ram_block1a175,
	ram_block1a55,
	ram_block1a79,
	ram_block1a7,
	ram_block1a31,
	ram_block1a104,
	ram_block1a128,
	ram_block1a152,
	ram_block1a176,
	ram_block1a56,
	ram_block1a80,
	ram_block1a8,
	ram_block1a32,
	ram_block1a105,
	ram_block1a129,
	ram_block1a153,
	ram_block1a177,
	ram_block1a57,
	ram_block1a81,
	ram_block1a9,
	ram_block1a33,
	ram_block1a106,
	ram_block1a130,
	ram_block1a154,
	ram_block1a178,
	ram_block1a58,
	ram_block1a82,
	ram_block1a10,
	ram_block1a34,
	ram_block1a107,
	ram_block1a131,
	ram_block1a155,
	ram_block1a179,
	ram_block1a59,
	ram_block1a83,
	ram_block1a11,
	ram_block1a35,
	ram_block1a108,
	ram_block1a132,
	ram_block1a156,
	ram_block1a180,
	ram_block1a60,
	ram_block1a84,
	ram_block1a12,
	ram_block1a36,
	ram_block1a109,
	ram_block1a133,
	ram_block1a157,
	ram_block1a181,
	ram_block1a61,
	ram_block1a85,
	ram_block1a13,
	ram_block1a37,
	ram_block1a110,
	ram_block1a134,
	ram_block1a158,
	ram_block1a182,
	ram_block1a62,
	ram_block1a86,
	ram_block1a14,
	ram_block1a38,
	ram_block1a111,
	ram_block1a135,
	ram_block1a159,
	ram_block1a183,
	ram_block1a63,
	ram_block1a87,
	ram_block1a15,
	ram_block1a39,
	ram_block1a112,
	ram_block1a136,
	ram_block1a160,
	ram_block1a184,
	ram_block1a64,
	ram_block1a88,
	ram_block1a16,
	ram_block1a40,
	ram_block1a113,
	ram_block1a137,
	ram_block1a161,
	ram_block1a185,
	ram_block1a65,
	ram_block1a89,
	ram_block1a17,
	ram_block1a41,
	ram_block1a114,
	ram_block1a138,
	ram_block1a162,
	ram_block1a186,
	ram_block1a66,
	ram_block1a90,
	ram_block1a18,
	ram_block1a42,
	ram_block1a115,
	ram_block1a139,
	ram_block1a163,
	ram_block1a187,
	ram_block1a67,
	ram_block1a91,
	ram_block1a19,
	ram_block1a43,
	ram_block1a116,
	ram_block1a140,
	ram_block1a164,
	ram_block1a188,
	ram_block1a68,
	ram_block1a92,
	ram_block1a20,
	ram_block1a44,
	ram_block1a117,
	ram_block1a141,
	ram_block1a165,
	ram_block1a189,
	ram_block1a69,
	ram_block1a93,
	ram_block1a21,
	ram_block1a45,
	ram_block1a118,
	ram_block1a142,
	ram_block1a166,
	ram_block1a190,
	ram_block1a70,
	ram_block1a94,
	ram_block1a22,
	ram_block1a46,
	ram_block1a119,
	ram_block1a143,
	ram_block1a167,
	ram_block1a191,
	ram_block1a71,
	ram_block1a95,
	ram_block1a23,
	ram_block1a47,
	out_address_reg_a_2,
	out_address_reg_a_0,
	out_address_reg_a_1,
	data_out_121,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
output 	data_out_8;
output 	data_out_9;
output 	data_out_10;
output 	data_out_11;
output 	data_out_12;
output 	data_out_13;
output 	data_out_14;
output 	data_out_15;
output 	data_out_16;
output 	data_out_17;
output 	data_out_18;
output 	data_out_19;
output 	data_out_20;
output 	data_out_21;
output 	data_out_22;
output 	data_out_23;
input 	ram_block1a96;
input 	ram_block1a120;
input 	ram_block1a144;
input 	ram_block1a168;
input 	ram_block1a48;
input 	ram_block1a72;
input 	ram_block1a0;
input 	ram_block1a24;
input 	ram_block1a97;
input 	ram_block1a121;
input 	ram_block1a145;
input 	ram_block1a169;
input 	ram_block1a49;
input 	ram_block1a73;
input 	ram_block1a1;
input 	ram_block1a25;
input 	ram_block1a98;
input 	ram_block1a122;
input 	ram_block1a146;
input 	ram_block1a170;
input 	ram_block1a50;
input 	ram_block1a74;
input 	ram_block1a2;
input 	ram_block1a26;
input 	ram_block1a99;
input 	ram_block1a123;
input 	ram_block1a147;
input 	ram_block1a171;
input 	ram_block1a51;
input 	ram_block1a75;
input 	ram_block1a3;
input 	ram_block1a27;
input 	ram_block1a100;
input 	ram_block1a124;
input 	ram_block1a148;
input 	ram_block1a172;
input 	ram_block1a52;
input 	ram_block1a76;
input 	ram_block1a4;
input 	ram_block1a28;
input 	ram_block1a101;
input 	ram_block1a125;
input 	ram_block1a149;
input 	ram_block1a173;
input 	ram_block1a53;
input 	ram_block1a77;
input 	ram_block1a5;
input 	ram_block1a29;
input 	ram_block1a102;
input 	ram_block1a126;
input 	ram_block1a150;
input 	ram_block1a174;
input 	ram_block1a54;
input 	ram_block1a78;
input 	ram_block1a6;
input 	ram_block1a30;
input 	ram_block1a103;
input 	ram_block1a127;
input 	ram_block1a151;
input 	ram_block1a175;
input 	ram_block1a55;
input 	ram_block1a79;
input 	ram_block1a7;
input 	ram_block1a31;
input 	ram_block1a104;
input 	ram_block1a128;
input 	ram_block1a152;
input 	ram_block1a176;
input 	ram_block1a56;
input 	ram_block1a80;
input 	ram_block1a8;
input 	ram_block1a32;
input 	ram_block1a105;
input 	ram_block1a129;
input 	ram_block1a153;
input 	ram_block1a177;
input 	ram_block1a57;
input 	ram_block1a81;
input 	ram_block1a9;
input 	ram_block1a33;
input 	ram_block1a106;
input 	ram_block1a130;
input 	ram_block1a154;
input 	ram_block1a178;
input 	ram_block1a58;
input 	ram_block1a82;
input 	ram_block1a10;
input 	ram_block1a34;
input 	ram_block1a107;
input 	ram_block1a131;
input 	ram_block1a155;
input 	ram_block1a179;
input 	ram_block1a59;
input 	ram_block1a83;
input 	ram_block1a11;
input 	ram_block1a35;
input 	ram_block1a108;
input 	ram_block1a132;
input 	ram_block1a156;
input 	ram_block1a180;
input 	ram_block1a60;
input 	ram_block1a84;
input 	ram_block1a12;
input 	ram_block1a36;
input 	ram_block1a109;
input 	ram_block1a133;
input 	ram_block1a157;
input 	ram_block1a181;
input 	ram_block1a61;
input 	ram_block1a85;
input 	ram_block1a13;
input 	ram_block1a37;
input 	ram_block1a110;
input 	ram_block1a134;
input 	ram_block1a158;
input 	ram_block1a182;
input 	ram_block1a62;
input 	ram_block1a86;
input 	ram_block1a14;
input 	ram_block1a38;
input 	ram_block1a111;
input 	ram_block1a135;
input 	ram_block1a159;
input 	ram_block1a183;
input 	ram_block1a63;
input 	ram_block1a87;
input 	ram_block1a15;
input 	ram_block1a39;
input 	ram_block1a112;
input 	ram_block1a136;
input 	ram_block1a160;
input 	ram_block1a184;
input 	ram_block1a64;
input 	ram_block1a88;
input 	ram_block1a16;
input 	ram_block1a40;
input 	ram_block1a113;
input 	ram_block1a137;
input 	ram_block1a161;
input 	ram_block1a185;
input 	ram_block1a65;
input 	ram_block1a89;
input 	ram_block1a17;
input 	ram_block1a41;
input 	ram_block1a114;
input 	ram_block1a138;
input 	ram_block1a162;
input 	ram_block1a186;
input 	ram_block1a66;
input 	ram_block1a90;
input 	ram_block1a18;
input 	ram_block1a42;
input 	ram_block1a115;
input 	ram_block1a139;
input 	ram_block1a163;
input 	ram_block1a187;
input 	ram_block1a67;
input 	ram_block1a91;
input 	ram_block1a19;
input 	ram_block1a43;
input 	ram_block1a116;
input 	ram_block1a140;
input 	ram_block1a164;
input 	ram_block1a188;
input 	ram_block1a68;
input 	ram_block1a92;
input 	ram_block1a20;
input 	ram_block1a44;
input 	ram_block1a117;
input 	ram_block1a141;
input 	ram_block1a165;
input 	ram_block1a189;
input 	ram_block1a69;
input 	ram_block1a93;
input 	ram_block1a21;
input 	ram_block1a45;
input 	ram_block1a118;
input 	ram_block1a142;
input 	ram_block1a166;
input 	ram_block1a190;
input 	ram_block1a70;
input 	ram_block1a94;
input 	ram_block1a22;
input 	ram_block1a46;
input 	ram_block1a119;
input 	ram_block1a143;
input 	ram_block1a167;
input 	ram_block1a191;
input 	ram_block1a71;
input 	ram_block1a95;
input 	ram_block1a23;
input 	ram_block1a47;
input 	out_address_reg_a_2;
input 	out_address_reg_a_0;
input 	out_address_reg_a_1;
output 	data_out_121;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out~0_combout ;
wire \data_out~1_combout ;
wire \data_out~2_combout ;
wire \data_out~4_combout ;
wire \data_out~5_combout ;
wire \data_out~6_combout ;
wire \data_out~7_combout ;
wire \data_out~8_combout ;
wire \data_out~9_combout ;
wire \data_out~10_combout ;
wire \data_out~11_combout ;
wire \data_out~12_combout ;
wire \data_out~13_combout ;
wire \data_out~14_combout ;
wire \data_out~15_combout ;
wire \data_out~16_combout ;
wire \data_out~17_combout ;
wire \data_out~18_combout ;
wire \data_out~19_combout ;
wire \data_out~20_combout ;
wire \data_out~21_combout ;
wire \data_out~22_combout ;
wire \data_out~23_combout ;
wire \data_out~24_combout ;
wire \data_out~25_combout ;
wire \data_out~26_combout ;
wire \data_out~27_combout ;
wire \data_out~28_combout ;
wire \data_out~29_combout ;
wire \data_out~30_combout ;
wire \data_out~31_combout ;
wire \data_out~32_combout ;
wire \data_out~33_combout ;
wire \data_out~34_combout ;
wire \data_out~35_combout ;
wire \data_out~36_combout ;
wire \data_out~37_combout ;
wire \data_out~38_combout ;
wire \data_out~39_combout ;
wire \data_out~40_combout ;
wire \data_out~41_combout ;
wire \data_out~42_combout ;
wire \data_out~43_combout ;
wire \data_out~44_combout ;
wire \data_out~45_combout ;
wire \data_out~46_combout ;
wire \data_out~47_combout ;
wire \data_out~48_combout ;
wire \data_out~49_combout ;
wire \data_out~50_combout ;
wire \data_out~51_combout ;
wire \data_out~52_combout ;
wire \data_out~53_combout ;
wire \data_out~54_combout ;
wire \data_out~55_combout ;
wire \data_out~56_combout ;
wire \data_out~57_combout ;
wire \data_out~58_combout ;
wire \data_out~59_combout ;
wire \data_out~60_combout ;
wire \data_out~61_combout ;
wire \data_out~62_combout ;
wire \data_out~63_combout ;
wire \data_out~64_combout ;
wire \data_out~65_combout ;
wire \data_out~66_combout ;
wire \data_out~67_combout ;
wire \data_out~68_combout ;
wire \data_out~69_combout ;
wire \data_out~70_combout ;
wire \data_out~71_combout ;
wire \data_out~72_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(\data_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(\data_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(\data_out~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(\data_out~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(\data_out~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(\data_out~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(\data_out~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(\data_out~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk),
	.d(\data_out~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

dffeas \data_out[9] (
	.clk(clk),
	.d(\data_out~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_9),
	.prn(vcc));
defparam \data_out[9] .is_wysiwyg = "true";
defparam \data_out[9] .power_up = "low";

dffeas \data_out[10] (
	.clk(clk),
	.d(\data_out~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_10),
	.prn(vcc));
defparam \data_out[10] .is_wysiwyg = "true";
defparam \data_out[10] .power_up = "low";

dffeas \data_out[11] (
	.clk(clk),
	.d(\data_out~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_11),
	.prn(vcc));
defparam \data_out[11] .is_wysiwyg = "true";
defparam \data_out[11] .power_up = "low";

dffeas \data_out[12] (
	.clk(clk),
	.d(\data_out~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_12),
	.prn(vcc));
defparam \data_out[12] .is_wysiwyg = "true";
defparam \data_out[12] .power_up = "low";

dffeas \data_out[13] (
	.clk(clk),
	.d(\data_out~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_13),
	.prn(vcc));
defparam \data_out[13] .is_wysiwyg = "true";
defparam \data_out[13] .power_up = "low";

dffeas \data_out[14] (
	.clk(clk),
	.d(\data_out~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_14),
	.prn(vcc));
defparam \data_out[14] .is_wysiwyg = "true";
defparam \data_out[14] .power_up = "low";

dffeas \data_out[15] (
	.clk(clk),
	.d(\data_out~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_15),
	.prn(vcc));
defparam \data_out[15] .is_wysiwyg = "true";
defparam \data_out[15] .power_up = "low";

dffeas \data_out[16] (
	.clk(clk),
	.d(\data_out~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_16),
	.prn(vcc));
defparam \data_out[16] .is_wysiwyg = "true";
defparam \data_out[16] .power_up = "low";

dffeas \data_out[17] (
	.clk(clk),
	.d(\data_out~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_17),
	.prn(vcc));
defparam \data_out[17] .is_wysiwyg = "true";
defparam \data_out[17] .power_up = "low";

dffeas \data_out[18] (
	.clk(clk),
	.d(\data_out~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_18),
	.prn(vcc));
defparam \data_out[18] .is_wysiwyg = "true";
defparam \data_out[18] .power_up = "low";

dffeas \data_out[19] (
	.clk(clk),
	.d(\data_out~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_19),
	.prn(vcc));
defparam \data_out[19] .is_wysiwyg = "true";
defparam \data_out[19] .power_up = "low";

dffeas \data_out[20] (
	.clk(clk),
	.d(\data_out~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_20),
	.prn(vcc));
defparam \data_out[20] .is_wysiwyg = "true";
defparam \data_out[20] .power_up = "low";

dffeas \data_out[21] (
	.clk(clk),
	.d(\data_out~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_21),
	.prn(vcc));
defparam \data_out[21] .is_wysiwyg = "true";
defparam \data_out[21] .power_up = "low";

dffeas \data_out[22] (
	.clk(clk),
	.d(\data_out~69_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_22),
	.prn(vcc));
defparam \data_out[22] .is_wysiwyg = "true";
defparam \data_out[22] .power_up = "low";

dffeas \data_out[23] (
	.clk(clk),
	.d(\data_out~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_121),
	.q(data_out_23),
	.prn(vcc));
defparam \data_out[23] .is_wysiwyg = "true";
defparam \data_out[23] .power_up = "low";

cyclonev_lcell_comb \data_out[12]~3 (
	.dataa(!reset_n),
	.datab(!clken),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(data_out_121),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out[12]~3 .extended_lut = "off";
defparam \data_out[12]~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \data_out[12]~3 .shared_arith = "off";

cyclonev_lcell_comb \data_out~0 (
	.dataa(!ram_block1a96),
	.datab(!ram_block1a120),
	.datac(!ram_block1a144),
	.datad(!ram_block1a168),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~0 .extended_lut = "off";
defparam \data_out~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~0 .shared_arith = "off";

cyclonev_lcell_comb \data_out~1 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a48),
	.datad(!ram_block1a72),
	.datae(!ram_block1a0),
	.dataf(!ram_block1a24),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~1 .extended_lut = "off";
defparam \data_out~1 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~1 .shared_arith = "off";

cyclonev_lcell_comb \data_out~2 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~0_combout ),
	.datac(!\data_out~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~2 .extended_lut = "off";
defparam \data_out~2 .lut_mask = 64'h2727272727272727;
defparam \data_out~2 .shared_arith = "off";

cyclonev_lcell_comb \data_out~4 (
	.dataa(!ram_block1a97),
	.datab(!ram_block1a121),
	.datac(!ram_block1a145),
	.datad(!ram_block1a169),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~4 .extended_lut = "off";
defparam \data_out~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~4 .shared_arith = "off";

cyclonev_lcell_comb \data_out~5 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a49),
	.datad(!ram_block1a73),
	.datae(!ram_block1a1),
	.dataf(!ram_block1a25),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~5 .extended_lut = "off";
defparam \data_out~5 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~5 .shared_arith = "off";

cyclonev_lcell_comb \data_out~6 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~4_combout ),
	.datac(!\data_out~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~6 .extended_lut = "off";
defparam \data_out~6 .lut_mask = 64'h2727272727272727;
defparam \data_out~6 .shared_arith = "off";

cyclonev_lcell_comb \data_out~7 (
	.dataa(!ram_block1a98),
	.datab(!ram_block1a122),
	.datac(!ram_block1a146),
	.datad(!ram_block1a170),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~7 .extended_lut = "off";
defparam \data_out~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~7 .shared_arith = "off";

cyclonev_lcell_comb \data_out~8 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a50),
	.datad(!ram_block1a74),
	.datae(!ram_block1a2),
	.dataf(!ram_block1a26),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~8 .extended_lut = "off";
defparam \data_out~8 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~8 .shared_arith = "off";

cyclonev_lcell_comb \data_out~9 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~7_combout ),
	.datac(!\data_out~8_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~9 .extended_lut = "off";
defparam \data_out~9 .lut_mask = 64'h2727272727272727;
defparam \data_out~9 .shared_arith = "off";

cyclonev_lcell_comb \data_out~10 (
	.dataa(!ram_block1a99),
	.datab(!ram_block1a123),
	.datac(!ram_block1a147),
	.datad(!ram_block1a171),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~10 .extended_lut = "off";
defparam \data_out~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~10 .shared_arith = "off";

cyclonev_lcell_comb \data_out~11 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a51),
	.datad(!ram_block1a75),
	.datae(!ram_block1a3),
	.dataf(!ram_block1a27),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~11 .extended_lut = "off";
defparam \data_out~11 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~11 .shared_arith = "off";

cyclonev_lcell_comb \data_out~12 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~10_combout ),
	.datac(!\data_out~11_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~12 .extended_lut = "off";
defparam \data_out~12 .lut_mask = 64'h2727272727272727;
defparam \data_out~12 .shared_arith = "off";

cyclonev_lcell_comb \data_out~13 (
	.dataa(!ram_block1a100),
	.datab(!ram_block1a124),
	.datac(!ram_block1a148),
	.datad(!ram_block1a172),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~13 .extended_lut = "off";
defparam \data_out~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~13 .shared_arith = "off";

cyclonev_lcell_comb \data_out~14 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a52),
	.datad(!ram_block1a76),
	.datae(!ram_block1a4),
	.dataf(!ram_block1a28),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~14 .extended_lut = "off";
defparam \data_out~14 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~14 .shared_arith = "off";

cyclonev_lcell_comb \data_out~15 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~13_combout ),
	.datac(!\data_out~14_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~15 .extended_lut = "off";
defparam \data_out~15 .lut_mask = 64'h2727272727272727;
defparam \data_out~15 .shared_arith = "off";

cyclonev_lcell_comb \data_out~16 (
	.dataa(!ram_block1a101),
	.datab(!ram_block1a125),
	.datac(!ram_block1a149),
	.datad(!ram_block1a173),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~16 .extended_lut = "off";
defparam \data_out~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~16 .shared_arith = "off";

cyclonev_lcell_comb \data_out~17 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a53),
	.datad(!ram_block1a77),
	.datae(!ram_block1a5),
	.dataf(!ram_block1a29),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~17 .extended_lut = "off";
defparam \data_out~17 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~17 .shared_arith = "off";

cyclonev_lcell_comb \data_out~18 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~16_combout ),
	.datac(!\data_out~17_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~18 .extended_lut = "off";
defparam \data_out~18 .lut_mask = 64'h2727272727272727;
defparam \data_out~18 .shared_arith = "off";

cyclonev_lcell_comb \data_out~19 (
	.dataa(!ram_block1a102),
	.datab(!ram_block1a126),
	.datac(!ram_block1a150),
	.datad(!ram_block1a174),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~19 .extended_lut = "off";
defparam \data_out~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~19 .shared_arith = "off";

cyclonev_lcell_comb \data_out~20 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a54),
	.datad(!ram_block1a78),
	.datae(!ram_block1a6),
	.dataf(!ram_block1a30),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~20 .extended_lut = "off";
defparam \data_out~20 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~20 .shared_arith = "off";

cyclonev_lcell_comb \data_out~21 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~19_combout ),
	.datac(!\data_out~20_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~21 .extended_lut = "off";
defparam \data_out~21 .lut_mask = 64'h2727272727272727;
defparam \data_out~21 .shared_arith = "off";

cyclonev_lcell_comb \data_out~22 (
	.dataa(!ram_block1a103),
	.datab(!ram_block1a127),
	.datac(!ram_block1a151),
	.datad(!ram_block1a175),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~22 .extended_lut = "off";
defparam \data_out~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~22 .shared_arith = "off";

cyclonev_lcell_comb \data_out~23 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a55),
	.datad(!ram_block1a79),
	.datae(!ram_block1a7),
	.dataf(!ram_block1a31),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~23 .extended_lut = "off";
defparam \data_out~23 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~23 .shared_arith = "off";

cyclonev_lcell_comb \data_out~24 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~22_combout ),
	.datac(!\data_out~23_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~24 .extended_lut = "off";
defparam \data_out~24 .lut_mask = 64'h2727272727272727;
defparam \data_out~24 .shared_arith = "off";

cyclonev_lcell_comb \data_out~25 (
	.dataa(!ram_block1a104),
	.datab(!ram_block1a128),
	.datac(!ram_block1a152),
	.datad(!ram_block1a176),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~25 .extended_lut = "off";
defparam \data_out~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~25 .shared_arith = "off";

cyclonev_lcell_comb \data_out~26 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a56),
	.datad(!ram_block1a80),
	.datae(!ram_block1a8),
	.dataf(!ram_block1a32),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~26 .extended_lut = "off";
defparam \data_out~26 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~26 .shared_arith = "off";

cyclonev_lcell_comb \data_out~27 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~25_combout ),
	.datac(!\data_out~26_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~27 .extended_lut = "off";
defparam \data_out~27 .lut_mask = 64'h2727272727272727;
defparam \data_out~27 .shared_arith = "off";

cyclonev_lcell_comb \data_out~28 (
	.dataa(!ram_block1a105),
	.datab(!ram_block1a129),
	.datac(!ram_block1a153),
	.datad(!ram_block1a177),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~28 .extended_lut = "off";
defparam \data_out~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~28 .shared_arith = "off";

cyclonev_lcell_comb \data_out~29 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a57),
	.datad(!ram_block1a81),
	.datae(!ram_block1a9),
	.dataf(!ram_block1a33),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~29 .extended_lut = "off";
defparam \data_out~29 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~29 .shared_arith = "off";

cyclonev_lcell_comb \data_out~30 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~28_combout ),
	.datac(!\data_out~29_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~30 .extended_lut = "off";
defparam \data_out~30 .lut_mask = 64'h2727272727272727;
defparam \data_out~30 .shared_arith = "off";

cyclonev_lcell_comb \data_out~31 (
	.dataa(!ram_block1a106),
	.datab(!ram_block1a130),
	.datac(!ram_block1a154),
	.datad(!ram_block1a178),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~31 .extended_lut = "off";
defparam \data_out~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~31 .shared_arith = "off";

cyclonev_lcell_comb \data_out~32 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a58),
	.datad(!ram_block1a82),
	.datae(!ram_block1a10),
	.dataf(!ram_block1a34),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~32 .extended_lut = "off";
defparam \data_out~32 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~32 .shared_arith = "off";

cyclonev_lcell_comb \data_out~33 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~31_combout ),
	.datac(!\data_out~32_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~33 .extended_lut = "off";
defparam \data_out~33 .lut_mask = 64'h2727272727272727;
defparam \data_out~33 .shared_arith = "off";

cyclonev_lcell_comb \data_out~34 (
	.dataa(!ram_block1a107),
	.datab(!ram_block1a131),
	.datac(!ram_block1a155),
	.datad(!ram_block1a179),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~34 .extended_lut = "off";
defparam \data_out~34 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~34 .shared_arith = "off";

cyclonev_lcell_comb \data_out~35 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a59),
	.datad(!ram_block1a83),
	.datae(!ram_block1a11),
	.dataf(!ram_block1a35),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~35 .extended_lut = "off";
defparam \data_out~35 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~35 .shared_arith = "off";

cyclonev_lcell_comb \data_out~36 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~34_combout ),
	.datac(!\data_out~35_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~36 .extended_lut = "off";
defparam \data_out~36 .lut_mask = 64'h2727272727272727;
defparam \data_out~36 .shared_arith = "off";

cyclonev_lcell_comb \data_out~37 (
	.dataa(!ram_block1a108),
	.datab(!ram_block1a132),
	.datac(!ram_block1a156),
	.datad(!ram_block1a180),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~37 .extended_lut = "off";
defparam \data_out~37 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~37 .shared_arith = "off";

cyclonev_lcell_comb \data_out~38 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a60),
	.datad(!ram_block1a84),
	.datae(!ram_block1a12),
	.dataf(!ram_block1a36),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~38 .extended_lut = "off";
defparam \data_out~38 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~38 .shared_arith = "off";

cyclonev_lcell_comb \data_out~39 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~37_combout ),
	.datac(!\data_out~38_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~39 .extended_lut = "off";
defparam \data_out~39 .lut_mask = 64'h2727272727272727;
defparam \data_out~39 .shared_arith = "off";

cyclonev_lcell_comb \data_out~40 (
	.dataa(!ram_block1a109),
	.datab(!ram_block1a133),
	.datac(!ram_block1a157),
	.datad(!ram_block1a181),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~40 .extended_lut = "off";
defparam \data_out~40 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~40 .shared_arith = "off";

cyclonev_lcell_comb \data_out~41 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a61),
	.datad(!ram_block1a85),
	.datae(!ram_block1a13),
	.dataf(!ram_block1a37),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~41 .extended_lut = "off";
defparam \data_out~41 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~41 .shared_arith = "off";

cyclonev_lcell_comb \data_out~42 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~40_combout ),
	.datac(!\data_out~41_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~42 .extended_lut = "off";
defparam \data_out~42 .lut_mask = 64'h2727272727272727;
defparam \data_out~42 .shared_arith = "off";

cyclonev_lcell_comb \data_out~43 (
	.dataa(!ram_block1a110),
	.datab(!ram_block1a134),
	.datac(!ram_block1a158),
	.datad(!ram_block1a182),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~43 .extended_lut = "off";
defparam \data_out~43 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~43 .shared_arith = "off";

cyclonev_lcell_comb \data_out~44 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a62),
	.datad(!ram_block1a86),
	.datae(!ram_block1a14),
	.dataf(!ram_block1a38),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~44 .extended_lut = "off";
defparam \data_out~44 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~44 .shared_arith = "off";

cyclonev_lcell_comb \data_out~45 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~43_combout ),
	.datac(!\data_out~44_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~45 .extended_lut = "off";
defparam \data_out~45 .lut_mask = 64'h2727272727272727;
defparam \data_out~45 .shared_arith = "off";

cyclonev_lcell_comb \data_out~46 (
	.dataa(!ram_block1a111),
	.datab(!ram_block1a135),
	.datac(!ram_block1a159),
	.datad(!ram_block1a183),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~46 .extended_lut = "off";
defparam \data_out~46 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~46 .shared_arith = "off";

cyclonev_lcell_comb \data_out~47 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a63),
	.datad(!ram_block1a87),
	.datae(!ram_block1a15),
	.dataf(!ram_block1a39),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~47 .extended_lut = "off";
defparam \data_out~47 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~47 .shared_arith = "off";

cyclonev_lcell_comb \data_out~48 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~46_combout ),
	.datac(!\data_out~47_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~48 .extended_lut = "off";
defparam \data_out~48 .lut_mask = 64'h2727272727272727;
defparam \data_out~48 .shared_arith = "off";

cyclonev_lcell_comb \data_out~49 (
	.dataa(!ram_block1a112),
	.datab(!ram_block1a136),
	.datac(!ram_block1a160),
	.datad(!ram_block1a184),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~49 .extended_lut = "off";
defparam \data_out~49 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~49 .shared_arith = "off";

cyclonev_lcell_comb \data_out~50 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a64),
	.datad(!ram_block1a88),
	.datae(!ram_block1a16),
	.dataf(!ram_block1a40),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~50 .extended_lut = "off";
defparam \data_out~50 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~50 .shared_arith = "off";

cyclonev_lcell_comb \data_out~51 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~49_combout ),
	.datac(!\data_out~50_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~51 .extended_lut = "off";
defparam \data_out~51 .lut_mask = 64'h2727272727272727;
defparam \data_out~51 .shared_arith = "off";

cyclonev_lcell_comb \data_out~52 (
	.dataa(!ram_block1a113),
	.datab(!ram_block1a137),
	.datac(!ram_block1a161),
	.datad(!ram_block1a185),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~52 .extended_lut = "off";
defparam \data_out~52 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~52 .shared_arith = "off";

cyclonev_lcell_comb \data_out~53 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a65),
	.datad(!ram_block1a89),
	.datae(!ram_block1a17),
	.dataf(!ram_block1a41),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~53 .extended_lut = "off";
defparam \data_out~53 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~53 .shared_arith = "off";

cyclonev_lcell_comb \data_out~54 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~52_combout ),
	.datac(!\data_out~53_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~54 .extended_lut = "off";
defparam \data_out~54 .lut_mask = 64'h2727272727272727;
defparam \data_out~54 .shared_arith = "off";

cyclonev_lcell_comb \data_out~55 (
	.dataa(!ram_block1a114),
	.datab(!ram_block1a138),
	.datac(!ram_block1a162),
	.datad(!ram_block1a186),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~55 .extended_lut = "off";
defparam \data_out~55 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~55 .shared_arith = "off";

cyclonev_lcell_comb \data_out~56 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a66),
	.datad(!ram_block1a90),
	.datae(!ram_block1a18),
	.dataf(!ram_block1a42),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~56 .extended_lut = "off";
defparam \data_out~56 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~56 .shared_arith = "off";

cyclonev_lcell_comb \data_out~57 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~55_combout ),
	.datac(!\data_out~56_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~57 .extended_lut = "off";
defparam \data_out~57 .lut_mask = 64'h2727272727272727;
defparam \data_out~57 .shared_arith = "off";

cyclonev_lcell_comb \data_out~58 (
	.dataa(!ram_block1a115),
	.datab(!ram_block1a139),
	.datac(!ram_block1a163),
	.datad(!ram_block1a187),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~58 .extended_lut = "off";
defparam \data_out~58 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~58 .shared_arith = "off";

cyclonev_lcell_comb \data_out~59 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a67),
	.datad(!ram_block1a91),
	.datae(!ram_block1a19),
	.dataf(!ram_block1a43),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~59 .extended_lut = "off";
defparam \data_out~59 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~59 .shared_arith = "off";

cyclonev_lcell_comb \data_out~60 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~58_combout ),
	.datac(!\data_out~59_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~60 .extended_lut = "off";
defparam \data_out~60 .lut_mask = 64'h2727272727272727;
defparam \data_out~60 .shared_arith = "off";

cyclonev_lcell_comb \data_out~61 (
	.dataa(!ram_block1a116),
	.datab(!ram_block1a140),
	.datac(!ram_block1a164),
	.datad(!ram_block1a188),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~61 .extended_lut = "off";
defparam \data_out~61 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~61 .shared_arith = "off";

cyclonev_lcell_comb \data_out~62 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a68),
	.datad(!ram_block1a92),
	.datae(!ram_block1a20),
	.dataf(!ram_block1a44),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~62 .extended_lut = "off";
defparam \data_out~62 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~62 .shared_arith = "off";

cyclonev_lcell_comb \data_out~63 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~61_combout ),
	.datac(!\data_out~62_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~63 .extended_lut = "off";
defparam \data_out~63 .lut_mask = 64'h2727272727272727;
defparam \data_out~63 .shared_arith = "off";

cyclonev_lcell_comb \data_out~64 (
	.dataa(!ram_block1a117),
	.datab(!ram_block1a141),
	.datac(!ram_block1a165),
	.datad(!ram_block1a189),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~64 .extended_lut = "off";
defparam \data_out~64 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~64 .shared_arith = "off";

cyclonev_lcell_comb \data_out~65 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a69),
	.datad(!ram_block1a93),
	.datae(!ram_block1a21),
	.dataf(!ram_block1a45),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~65 .extended_lut = "off";
defparam \data_out~65 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~65 .shared_arith = "off";

cyclonev_lcell_comb \data_out~66 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~64_combout ),
	.datac(!\data_out~65_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~66 .extended_lut = "off";
defparam \data_out~66 .lut_mask = 64'h2727272727272727;
defparam \data_out~66 .shared_arith = "off";

cyclonev_lcell_comb \data_out~67 (
	.dataa(!ram_block1a118),
	.datab(!ram_block1a142),
	.datac(!ram_block1a166),
	.datad(!ram_block1a190),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~67 .extended_lut = "off";
defparam \data_out~67 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~67 .shared_arith = "off";

cyclonev_lcell_comb \data_out~68 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a70),
	.datad(!ram_block1a94),
	.datae(!ram_block1a22),
	.dataf(!ram_block1a46),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~68 .extended_lut = "off";
defparam \data_out~68 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~68 .shared_arith = "off";

cyclonev_lcell_comb \data_out~69 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~67_combout ),
	.datac(!\data_out~68_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~69 .extended_lut = "off";
defparam \data_out~69 .lut_mask = 64'h2727272727272727;
defparam \data_out~69 .shared_arith = "off";

cyclonev_lcell_comb \data_out~70 (
	.dataa(!ram_block1a119),
	.datab(!ram_block1a143),
	.datac(!ram_block1a167),
	.datad(!ram_block1a191),
	.datae(!out_address_reg_a_0),
	.dataf(!out_address_reg_a_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~70 .extended_lut = "off";
defparam \data_out~70 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \data_out~70 .shared_arith = "off";

cyclonev_lcell_comb \data_out~71 (
	.dataa(!out_address_reg_a_0),
	.datab(!out_address_reg_a_1),
	.datac(!ram_block1a71),
	.datad(!ram_block1a95),
	.datae(!ram_block1a23),
	.dataf(!ram_block1a47),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~71_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~71 .extended_lut = "off";
defparam \data_out~71 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \data_out~71 .shared_arith = "off";

cyclonev_lcell_comb \data_out~72 (
	.dataa(!out_address_reg_a_2),
	.datab(!\data_out~70_combout ),
	.datac(!\data_out~71_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_out~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_out~72 .extended_lut = "off";
defparam \data_out~72 .lut_mask = 64'h2727272727272727;
defparam \data_out~72 .shared_arith = "off";

endmodule

module sine_asj_nco_pxx (
	dxxpdo_5,
	dxxpdo_6,
	dxxpdo_7,
	dxxpdo_8,
	dxxpdo_9,
	dxxpdo_10,
	dxxpdo_11,
	dxxpdo_12,
	dxxpdo_13,
	dxxpdo_14,
	dxxpdo_15,
	dxxpdo_16,
	dxxpdo_17,
	dxxpdo_20,
	dxxpdo_18,
	dxxpdo_19,
	data_out_12,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_15,
	pipeline_dffe_13,
	pipeline_dffe_14,
	clk,
	reset_n,
	clken,
	phase_mod_i_0,
	phase_mod_i_1,
	phase_mod_i_2,
	phase_mod_i_3,
	phase_mod_i_4,
	phase_mod_i_5,
	phase_mod_i_6,
	phase_mod_i_7,
	phase_mod_i_8,
	phase_mod_i_9,
	phase_mod_i_10,
	phase_mod_i_11,
	phase_mod_i_12,
	phase_mod_i_15,
	phase_mod_i_13,
	phase_mod_i_14)/* synthesis synthesis_greybox=1 */;
input 	dxxpdo_5;
input 	dxxpdo_6;
input 	dxxpdo_7;
input 	dxxpdo_8;
input 	dxxpdo_9;
input 	dxxpdo_10;
input 	dxxpdo_11;
input 	dxxpdo_12;
input 	dxxpdo_13;
input 	dxxpdo_14;
input 	dxxpdo_15;
input 	dxxpdo_16;
input 	dxxpdo_17;
input 	dxxpdo_20;
input 	dxxpdo_18;
input 	dxxpdo_19;
input 	data_out_12;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_15;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	clk;
input 	reset_n;
input 	clken;
input 	phase_mod_i_0;
input 	phase_mod_i_1;
input 	phase_mod_i_2;
input 	phase_mod_i_3;
input 	phase_mod_i_4;
input 	phase_mod_i_5;
input 	phase_mod_i_6;
input 	phase_mod_i_7;
input 	phase_mod_i_8;
input 	phase_mod_i_9;
input 	phase_mod_i_10;
input 	phase_mod_i_11;
input 	phase_mod_i_12;
input 	phase_mod_i_15;
input 	phase_mod_i_13;
input 	phase_mod_i_14;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \phi_mod_int_reg[3][0]~q ;
wire \phi_mod_int_reg[3][1]~q ;
wire \phi_mod_int_reg[3][2]~q ;
wire \phi_mod_int_reg[3][3]~q ;
wire \phi_mod_int_reg[3][4]~q ;
wire \phi_mod_int_reg[3][5]~q ;
wire \phi_mod_int_reg[3][6]~q ;
wire \phi_mod_int_reg[3][7]~q ;
wire \phi_mod_int_reg[3][8]~q ;
wire \phi_mod_int_reg[3][9]~q ;
wire \phi_mod_int_reg[3][10]~q ;
wire \phi_mod_int_reg[3][11]~q ;
wire \phi_mod_int_reg[3][12]~q ;
wire \phi_mod_int_reg[3][15]~q ;
wire \phi_mod_int_reg[2][0]~q ;
wire \phi_mod_int_reg[2][1]~q ;
wire \phi_mod_int_reg[2][2]~q ;
wire \phi_mod_int_reg[2][3]~q ;
wire \phi_mod_int_reg[2][4]~q ;
wire \phi_mod_int_reg[2][5]~q ;
wire \phi_mod_int_reg[2][6]~q ;
wire \phi_mod_int_reg[2][7]~q ;
wire \phi_mod_int_reg[2][8]~q ;
wire \phi_mod_int_reg[2][9]~q ;
wire \phi_mod_int_reg[2][10]~q ;
wire \phi_mod_int_reg[2][11]~q ;
wire \phi_mod_int_reg[2][12]~q ;
wire \phi_mod_int_reg[3][13]~q ;
wire \phi_mod_int_reg[3][14]~q ;
wire \phi_mod_int_reg[2][15]~q ;
wire \phi_mod_int_reg[1][0]~q ;
wire \phi_mod_int_reg[1][1]~q ;
wire \phi_mod_int_reg[1][2]~q ;
wire \phi_mod_int_reg[1][3]~q ;
wire \phi_mod_int_reg[1][4]~q ;
wire \phi_mod_int_reg[1][5]~q ;
wire \phi_mod_int_reg[1][6]~q ;
wire \phi_mod_int_reg[1][7]~q ;
wire \phi_mod_int_reg[1][8]~q ;
wire \phi_mod_int_reg[1][9]~q ;
wire \phi_mod_int_reg[1][10]~q ;
wire \phi_mod_int_reg[1][11]~q ;
wire \phi_mod_int_reg[1][12]~q ;
wire \phi_mod_int_reg[2][13]~q ;
wire \phi_mod_int_reg[2][14]~q ;
wire \phi_mod_int_reg[1][15]~q ;
wire \phi_mod_int_reg[0][0]~q ;
wire \phi_mod_int_reg[0][1]~q ;
wire \phi_mod_int_reg[0][2]~q ;
wire \phi_mod_int_reg[0][3]~q ;
wire \phi_mod_int_reg[0][4]~q ;
wire \phi_mod_int_reg[0][5]~q ;
wire \phi_mod_int_reg[0][6]~q ;
wire \phi_mod_int_reg[0][7]~q ;
wire \phi_mod_int_reg[0][8]~q ;
wire \phi_mod_int_reg[0][9]~q ;
wire \phi_mod_int_reg[0][10]~q ;
wire \phi_mod_int_reg[0][11]~q ;
wire \phi_mod_int_reg[0][12]~q ;
wire \phi_mod_int_reg[1][13]~q ;
wire \phi_mod_int_reg[1][14]~q ;
wire \phi_mod_int_reg[0][15]~q ;
wire \phi_mod_int_reg[0][13]~q ;
wire \phi_mod_int_reg[0][14]~q ;


sine_lpm_add_sub_3 acc(
	.dxxpdo_5(dxxpdo_5),
	.phi_mod_int_reg_0_3(\phi_mod_int_reg[3][0]~q ),
	.dxxpdo_6(dxxpdo_6),
	.phi_mod_int_reg_1_3(\phi_mod_int_reg[3][1]~q ),
	.dxxpdo_7(dxxpdo_7),
	.phi_mod_int_reg_2_3(\phi_mod_int_reg[3][2]~q ),
	.dxxpdo_8(dxxpdo_8),
	.phi_mod_int_reg_3_3(\phi_mod_int_reg[3][3]~q ),
	.dxxpdo_9(dxxpdo_9),
	.phi_mod_int_reg_4_3(\phi_mod_int_reg[3][4]~q ),
	.dxxpdo_10(dxxpdo_10),
	.phi_mod_int_reg_5_3(\phi_mod_int_reg[3][5]~q ),
	.dxxpdo_11(dxxpdo_11),
	.phi_mod_int_reg_6_3(\phi_mod_int_reg[3][6]~q ),
	.dxxpdo_12(dxxpdo_12),
	.phi_mod_int_reg_7_3(\phi_mod_int_reg[3][7]~q ),
	.dxxpdo_13(dxxpdo_13),
	.phi_mod_int_reg_8_3(\phi_mod_int_reg[3][8]~q ),
	.dxxpdo_14(dxxpdo_14),
	.phi_mod_int_reg_9_3(\phi_mod_int_reg[3][9]~q ),
	.dxxpdo_15(dxxpdo_15),
	.phi_mod_int_reg_10_3(\phi_mod_int_reg[3][10]~q ),
	.dxxpdo_16(dxxpdo_16),
	.phi_mod_int_reg_11_3(\phi_mod_int_reg[3][11]~q ),
	.dxxpdo_17(dxxpdo_17),
	.phi_mod_int_reg_12_3(\phi_mod_int_reg[3][12]~q ),
	.dxxpdo_20(dxxpdo_20),
	.phi_mod_int_reg_15_3(\phi_mod_int_reg[3][15]~q ),
	.phi_mod_int_reg_13_3(\phi_mod_int_reg[3][13]~q ),
	.dxxpdo_18(dxxpdo_18),
	.dxxpdo_19(dxxpdo_19),
	.phi_mod_int_reg_14_3(\phi_mod_int_reg[3][14]~q ),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \phi_mod_int_reg[3][0] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][0]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][0] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][0] .power_up = "low";

dffeas \phi_mod_int_reg[3][1] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][1]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][1] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][1] .power_up = "low";

dffeas \phi_mod_int_reg[3][2] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][2]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][2] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][2] .power_up = "low";

dffeas \phi_mod_int_reg[3][3] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][3]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][3] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][3] .power_up = "low";

dffeas \phi_mod_int_reg[3][4] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][4]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][4] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][4] .power_up = "low";

dffeas \phi_mod_int_reg[3][5] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][5]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][5] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][5] .power_up = "low";

dffeas \phi_mod_int_reg[3][6] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][6]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][6] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][6] .power_up = "low";

dffeas \phi_mod_int_reg[3][7] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][7]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][7] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][7] .power_up = "low";

dffeas \phi_mod_int_reg[3][8] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][8]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][8] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][8] .power_up = "low";

dffeas \phi_mod_int_reg[3][9] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][9]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][9] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][9] .power_up = "low";

dffeas \phi_mod_int_reg[3][10] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][10]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][10] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][10] .power_up = "low";

dffeas \phi_mod_int_reg[3][11] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][11]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][11] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][11] .power_up = "low";

dffeas \phi_mod_int_reg[3][12] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][12]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][12] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][12] .power_up = "low";

dffeas \phi_mod_int_reg[3][15] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][15]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][15] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][15] .power_up = "low";

dffeas \phi_mod_int_reg[2][0] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][0]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][0] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][0] .power_up = "low";

dffeas \phi_mod_int_reg[2][1] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][1]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][1] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][1] .power_up = "low";

dffeas \phi_mod_int_reg[2][2] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][2]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][2] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][2] .power_up = "low";

dffeas \phi_mod_int_reg[2][3] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][3]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][3] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][3] .power_up = "low";

dffeas \phi_mod_int_reg[2][4] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][4]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][4] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][4] .power_up = "low";

dffeas \phi_mod_int_reg[2][5] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][5]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][5] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][5] .power_up = "low";

dffeas \phi_mod_int_reg[2][6] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][6]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][6] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][6] .power_up = "low";

dffeas \phi_mod_int_reg[2][7] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][7]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][7] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][7] .power_up = "low";

dffeas \phi_mod_int_reg[2][8] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][8]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][8] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][8] .power_up = "low";

dffeas \phi_mod_int_reg[2][9] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][9]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][9] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][9] .power_up = "low";

dffeas \phi_mod_int_reg[2][10] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][10]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][10] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][10] .power_up = "low";

dffeas \phi_mod_int_reg[2][11] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][11]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][11] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][11] .power_up = "low";

dffeas \phi_mod_int_reg[2][12] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][12]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][12] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][12] .power_up = "low";

dffeas \phi_mod_int_reg[3][13] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][13]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][13] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][13] .power_up = "low";

dffeas \phi_mod_int_reg[3][14] (
	.clk(clk),
	.d(\phi_mod_int_reg[2][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[3][14]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[3][14] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[3][14] .power_up = "low";

dffeas \phi_mod_int_reg[2][15] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][15]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][15] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][15] .power_up = "low";

dffeas \phi_mod_int_reg[1][0] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][0]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][0] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][0] .power_up = "low";

dffeas \phi_mod_int_reg[1][1] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][1]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][1] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][1] .power_up = "low";

dffeas \phi_mod_int_reg[1][2] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][2]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][2] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][2] .power_up = "low";

dffeas \phi_mod_int_reg[1][3] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][3]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][3] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][3] .power_up = "low";

dffeas \phi_mod_int_reg[1][4] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][4]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][4] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][4] .power_up = "low";

dffeas \phi_mod_int_reg[1][5] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][5]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][5] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][5] .power_up = "low";

dffeas \phi_mod_int_reg[1][6] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][6]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][6] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][6] .power_up = "low";

dffeas \phi_mod_int_reg[1][7] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][7]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][7] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][7] .power_up = "low";

dffeas \phi_mod_int_reg[1][8] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][8]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][8] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][8] .power_up = "low";

dffeas \phi_mod_int_reg[1][9] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][9]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][9] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][9] .power_up = "low";

dffeas \phi_mod_int_reg[1][10] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][10]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][10] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][10] .power_up = "low";

dffeas \phi_mod_int_reg[1][11] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][11]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][11] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][11] .power_up = "low";

dffeas \phi_mod_int_reg[1][12] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][12]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][12] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][12] .power_up = "low";

dffeas \phi_mod_int_reg[2][13] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][13]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][13] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][13] .power_up = "low";

dffeas \phi_mod_int_reg[2][14] (
	.clk(clk),
	.d(\phi_mod_int_reg[1][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[2][14]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[2][14] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[2][14] .power_up = "low";

dffeas \phi_mod_int_reg[1][15] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][15]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][15] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][15] .power_up = "low";

dffeas \phi_mod_int_reg[0][0] (
	.clk(clk),
	.d(phase_mod_i_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][0]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][0] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][0] .power_up = "low";

dffeas \phi_mod_int_reg[0][1] (
	.clk(clk),
	.d(phase_mod_i_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][1]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][1] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][1] .power_up = "low";

dffeas \phi_mod_int_reg[0][2] (
	.clk(clk),
	.d(phase_mod_i_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][2]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][2] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][2] .power_up = "low";

dffeas \phi_mod_int_reg[0][3] (
	.clk(clk),
	.d(phase_mod_i_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][3]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][3] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][3] .power_up = "low";

dffeas \phi_mod_int_reg[0][4] (
	.clk(clk),
	.d(phase_mod_i_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][4]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][4] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][4] .power_up = "low";

dffeas \phi_mod_int_reg[0][5] (
	.clk(clk),
	.d(phase_mod_i_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][5]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][5] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][5] .power_up = "low";

dffeas \phi_mod_int_reg[0][6] (
	.clk(clk),
	.d(phase_mod_i_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][6]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][6] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][6] .power_up = "low";

dffeas \phi_mod_int_reg[0][7] (
	.clk(clk),
	.d(phase_mod_i_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][7]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][7] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][7] .power_up = "low";

dffeas \phi_mod_int_reg[0][8] (
	.clk(clk),
	.d(phase_mod_i_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][8]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][8] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][8] .power_up = "low";

dffeas \phi_mod_int_reg[0][9] (
	.clk(clk),
	.d(phase_mod_i_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][9]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][9] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][9] .power_up = "low";

dffeas \phi_mod_int_reg[0][10] (
	.clk(clk),
	.d(phase_mod_i_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][10]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][10] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][10] .power_up = "low";

dffeas \phi_mod_int_reg[0][11] (
	.clk(clk),
	.d(phase_mod_i_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][11]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][11] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][11] .power_up = "low";

dffeas \phi_mod_int_reg[0][12] (
	.clk(clk),
	.d(phase_mod_i_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][12]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][12] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][12] .power_up = "low";

dffeas \phi_mod_int_reg[1][13] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][13]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][13] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][13] .power_up = "low";

dffeas \phi_mod_int_reg[1][14] (
	.clk(clk),
	.d(\phi_mod_int_reg[0][14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[1][14]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[1][14] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[1][14] .power_up = "low";

dffeas \phi_mod_int_reg[0][15] (
	.clk(clk),
	.d(phase_mod_i_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][15]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][15] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][15] .power_up = "low";

dffeas \phi_mod_int_reg[0][13] (
	.clk(clk),
	.d(phase_mod_i_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][13]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][13] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][13] .power_up = "low";

dffeas \phi_mod_int_reg[0][14] (
	.clk(clk),
	.d(phase_mod_i_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(data_out_12),
	.q(\phi_mod_int_reg[0][14]~q ),
	.prn(vcc));
defparam \phi_mod_int_reg[0][14] .is_wysiwyg = "true";
defparam \phi_mod_int_reg[0][14] .power_up = "low";

endmodule

module sine_lpm_add_sub_3 (
	dxxpdo_5,
	phi_mod_int_reg_0_3,
	dxxpdo_6,
	phi_mod_int_reg_1_3,
	dxxpdo_7,
	phi_mod_int_reg_2_3,
	dxxpdo_8,
	phi_mod_int_reg_3_3,
	dxxpdo_9,
	phi_mod_int_reg_4_3,
	dxxpdo_10,
	phi_mod_int_reg_5_3,
	dxxpdo_11,
	phi_mod_int_reg_6_3,
	dxxpdo_12,
	phi_mod_int_reg_7_3,
	dxxpdo_13,
	phi_mod_int_reg_8_3,
	dxxpdo_14,
	phi_mod_int_reg_9_3,
	dxxpdo_15,
	phi_mod_int_reg_10_3,
	dxxpdo_16,
	phi_mod_int_reg_11_3,
	dxxpdo_17,
	phi_mod_int_reg_12_3,
	dxxpdo_20,
	phi_mod_int_reg_15_3,
	phi_mod_int_reg_13_3,
	dxxpdo_18,
	dxxpdo_19,
	phi_mod_int_reg_14_3,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_15,
	pipeline_dffe_13,
	pipeline_dffe_14,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	dxxpdo_5;
input 	phi_mod_int_reg_0_3;
input 	dxxpdo_6;
input 	phi_mod_int_reg_1_3;
input 	dxxpdo_7;
input 	phi_mod_int_reg_2_3;
input 	dxxpdo_8;
input 	phi_mod_int_reg_3_3;
input 	dxxpdo_9;
input 	phi_mod_int_reg_4_3;
input 	dxxpdo_10;
input 	phi_mod_int_reg_5_3;
input 	dxxpdo_11;
input 	phi_mod_int_reg_6_3;
input 	dxxpdo_12;
input 	phi_mod_int_reg_7_3;
input 	dxxpdo_13;
input 	phi_mod_int_reg_8_3;
input 	dxxpdo_14;
input 	phi_mod_int_reg_9_3;
input 	dxxpdo_15;
input 	phi_mod_int_reg_10_3;
input 	dxxpdo_16;
input 	phi_mod_int_reg_11_3;
input 	dxxpdo_17;
input 	phi_mod_int_reg_12_3;
input 	dxxpdo_20;
input 	phi_mod_int_reg_15_3;
input 	phi_mod_int_reg_13_3;
input 	dxxpdo_18;
input 	dxxpdo_19;
input 	phi_mod_int_reg_14_3;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_15;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



sine_add_sub_s0h auto_generated(
	.dxxpdo_5(dxxpdo_5),
	.phi_mod_int_reg_0_3(phi_mod_int_reg_0_3),
	.dxxpdo_6(dxxpdo_6),
	.phi_mod_int_reg_1_3(phi_mod_int_reg_1_3),
	.dxxpdo_7(dxxpdo_7),
	.phi_mod_int_reg_2_3(phi_mod_int_reg_2_3),
	.dxxpdo_8(dxxpdo_8),
	.phi_mod_int_reg_3_3(phi_mod_int_reg_3_3),
	.dxxpdo_9(dxxpdo_9),
	.phi_mod_int_reg_4_3(phi_mod_int_reg_4_3),
	.dxxpdo_10(dxxpdo_10),
	.phi_mod_int_reg_5_3(phi_mod_int_reg_5_3),
	.dxxpdo_11(dxxpdo_11),
	.phi_mod_int_reg_6_3(phi_mod_int_reg_6_3),
	.dxxpdo_12(dxxpdo_12),
	.phi_mod_int_reg_7_3(phi_mod_int_reg_7_3),
	.dxxpdo_13(dxxpdo_13),
	.phi_mod_int_reg_8_3(phi_mod_int_reg_8_3),
	.dxxpdo_14(dxxpdo_14),
	.phi_mod_int_reg_9_3(phi_mod_int_reg_9_3),
	.dxxpdo_15(dxxpdo_15),
	.phi_mod_int_reg_10_3(phi_mod_int_reg_10_3),
	.dxxpdo_16(dxxpdo_16),
	.phi_mod_int_reg_11_3(phi_mod_int_reg_11_3),
	.dxxpdo_17(dxxpdo_17),
	.phi_mod_int_reg_12_3(phi_mod_int_reg_12_3),
	.dxxpdo_20(dxxpdo_20),
	.phi_mod_int_reg_15_3(phi_mod_int_reg_15_3),
	.phi_mod_int_reg_13_3(phi_mod_int_reg_13_3),
	.dxxpdo_18(dxxpdo_18),
	.dxxpdo_19(dxxpdo_19),
	.phi_mod_int_reg_14_3(phi_mod_int_reg_14_3),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module sine_add_sub_s0h (
	dxxpdo_5,
	phi_mod_int_reg_0_3,
	dxxpdo_6,
	phi_mod_int_reg_1_3,
	dxxpdo_7,
	phi_mod_int_reg_2_3,
	dxxpdo_8,
	phi_mod_int_reg_3_3,
	dxxpdo_9,
	phi_mod_int_reg_4_3,
	dxxpdo_10,
	phi_mod_int_reg_5_3,
	dxxpdo_11,
	phi_mod_int_reg_6_3,
	dxxpdo_12,
	phi_mod_int_reg_7_3,
	dxxpdo_13,
	phi_mod_int_reg_8_3,
	dxxpdo_14,
	phi_mod_int_reg_9_3,
	dxxpdo_15,
	phi_mod_int_reg_10_3,
	dxxpdo_16,
	phi_mod_int_reg_11_3,
	dxxpdo_17,
	phi_mod_int_reg_12_3,
	dxxpdo_20,
	phi_mod_int_reg_15_3,
	phi_mod_int_reg_13_3,
	dxxpdo_18,
	dxxpdo_19,
	phi_mod_int_reg_14_3,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_15,
	pipeline_dffe_13,
	pipeline_dffe_14,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	dxxpdo_5;
input 	phi_mod_int_reg_0_3;
input 	dxxpdo_6;
input 	phi_mod_int_reg_1_3;
input 	dxxpdo_7;
input 	phi_mod_int_reg_2_3;
input 	dxxpdo_8;
input 	phi_mod_int_reg_3_3;
input 	dxxpdo_9;
input 	phi_mod_int_reg_4_3;
input 	dxxpdo_10;
input 	phi_mod_int_reg_5_3;
input 	dxxpdo_11;
input 	phi_mod_int_reg_6_3;
input 	dxxpdo_12;
input 	phi_mod_int_reg_7_3;
input 	dxxpdo_13;
input 	phi_mod_int_reg_8_3;
input 	dxxpdo_14;
input 	phi_mod_int_reg_9_3;
input 	dxxpdo_15;
input 	phi_mod_int_reg_10_3;
input 	dxxpdo_16;
input 	phi_mod_int_reg_11_3;
input 	dxxpdo_17;
input 	phi_mod_int_reg_12_3;
input 	dxxpdo_20;
input 	phi_mod_int_reg_15_3;
input 	phi_mod_int_reg_13_3;
input 	dxxpdo_18;
input 	dxxpdo_19;
input 	phi_mod_int_reg_14_3;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_15;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~6 ;
wire \op_1~9_sumout ;
wire \op_1~10 ;
wire \op_1~13_sumout ;
wire \op_1~14 ;
wire \op_1~17_sumout ;
wire \op_1~18 ;
wire \op_1~21_sumout ;
wire \op_1~22 ;
wire \op_1~25_sumout ;
wire \op_1~26 ;
wire \op_1~29_sumout ;
wire \op_1~30 ;
wire \op_1~33_sumout ;
wire \op_1~34 ;
wire \op_1~37_sumout ;
wire \op_1~38 ;
wire \op_1~41_sumout ;
wire \op_1~42 ;
wire \op_1~45_sumout ;
wire \op_1~46 ;
wire \op_1~49_sumout ;
wire \op_1~50 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;


dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_5),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_0_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_6),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_1_3),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_7),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_2_3),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_8),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_3_3),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_9),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_4_3),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_10),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_5_3),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_11),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_6_3),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_12),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_7_3),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_13),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_8_3),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_14),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_9_3),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_15),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_10_3),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_16),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_11_3),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_17),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_12_3),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

cyclonev_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_mod_int_reg_13_3),
	.datae(gnd),
	.dataf(!dxxpdo_18),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

cyclonev_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_19),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_14_3),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

cyclonev_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxpdo_20),
	.datae(gnd),
	.dataf(!phi_mod_int_reg_15_3),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

endmodule
