// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 15.1
// ALTERA_TIMESTAMP:Thu Oct 22 14:04:25 PDT 2015
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kp1V0dbROR7KsJXxzQn15KAp48kSWuI5jB5WQju65hkJshHNbLs5oNI/bytCVHxA
Zvk/lnSVWjw/EBcOiQc8st6V45BQKD0Ro5ThORogXcR4g554tQQX87PrhuLw8uhJ
GqnWdFJHExlKm/tFOMYysNVkJUAqIfm6ixkAyrHklSA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11456)
Q9+TUl50BFhAPZsegF0WIsphLMAfq0uyImF/Bw3KqsDwCLty54K5pkfLak7vBOYH
IYviCKvzrYjTbIUAFSz2ov22nJSGTYNGQhb3GTJXIguL6Ualy2G+qKVhK8s/2wQT
wMgZqugc7u0HMqFkKwrSGdzLgx2JJre8MY89LeOu971osQ003I3xacFhHUi4JktY
sFfo0s475Z295SaSgTEKFhUhFqTLsiD4h3kPKv6LoxcJGnF5mUatVHIK6Zl/5Q75
LRw07RQTVcUp2EMmDAPVtpB0NbwbWzViLpDASCc97akPxuhx6DAovDeofOLb2L0I
Ktw9W1TpweHhCfCxTHtObzqmtxmGFSXQBK6gK+k+6JtbPSo9RhCu6nmUlZTWBqeN
gxfY19WkfF+40apJ33QLUty3zxvRkxkKW7xZYu+CDjVN6RLpoiTXcRPhrI+nMDgA
mVtXWmh8LnEhcjjQLJyuN80fpgjwLJxP2RMWofyFxNi5Lye2qtuOzmo4BnBmZERO
polXUPV/h1LhBFPhzWh3JhXz9exveB+4T0mEeH9rU7kYkwzQ4Zvf11V3WcpXJyiS
iBUZbzqKOuqBh4+tnc8zGVdvKw/Wkn7XyC4VZ4ROc59vaFmZVJhMKv17aGbeFSA0
hxNwZiB3wxABc5R4lY6LFWE0uFFTRTDBJJYW4JaMHSulKpZesnnJkmnMTaTY/jcG
IoC8p2zZKxWO5UGC0QvGeg3lojjWKO/ve0Ak03tRuEOLgXXSdc/QM8a8txWPLff5
fQvNJ+vqcHLoc1j3P/cheqqnHBcruo2OYHxvyscjwjJrMFPEBDFLNtqyItDSCuKu
fg+p4QJdhK/5OHRD+oFbZxi4A1U0K9nA1AWcY8YNyXjIGPg6L0oHnFkMYHNJpKnB
VCiRRLSzsCHrjVIS1UF35Ef3JM0Dxi8nP11MbOgb7TgPKZmoysfMW6vohqwvZT2g
uyRhQImDgtgF+MvufKtz14eDpQGvX32GxyBQ1C8EEnzXUSvCvVLX0ssov7J7Zzbf
ygnDMy1R88Akn+F9pq6oP7TUN8Asrmg1j4bHq/aYmXyr17gY2QLJQSH6B8nFKkzE
X59i19GNmzAbAAJdWr5J9NmqJcu10D3kKupDs1qWIfCzHuC7QiNuS8j/+6d+4jN5
sJ7QDLqEb1/VyBjinGXo1alsT/vQ0NxaV9Zp/PsygZE4LahsHRXZLnDxIm3/Fptd
CVIMIKBw0CnTjSE7WVIKC4UcQDnbTjkrRRXrMRn0Br4x34pPEkqghnuT2q7TH1Mh
cwT9RfLTXTH4lTXrZpWs5HC36ILAXepTlp9wKzdvbTRR7PvcnUtOsHobOrGgrSUt
dRc+Z+rFHkXgEQfifwL9aGoFupGLk9J0P1LhBsi01N6I/gxNdUlpruUa1bosUEsO
qQbdf7aECM0/VVbBga4JSimzhsqokTOQ6wTYbysuRDcVTVgWl3jwHfS+xDXS8oK6
/oihfSEoNTrYGymmx8DjhqxeyjfzgfRGx9u0QBedXQSEAI7glgo+OSQUfZcwEZmQ
qHJDsTa/lBxYRe9uDjjBLNXVYm4kZCqt6hrRMEeFVazz11pkd5kokloX5RoEGHJY
UdK/rOB7fPPX5MHlYJ4ta9jPpF2cGpsntf+eK4TYpweqOxwv8gHT1yxAeMeD9wHr
mFCP2PABRAFSKToUXnErrf4evdnBFk+bwvhWOlusy0BYcglGi7kmDKPcOI2AU+hv
3jghyoMjTxlnb4XABEFRsqG7h/lrlFAcqhoP0VI/GQF+Ku8qjn8jAJfT4eOVAFer
hkl9fZQs3eyxDzu8XXXWom/dv2WoLUFFdE4xqDiJgZ+5CppbkBtyUcsm2JL2M1ar
wyuDKTzLB04ppL//4BgZvKGwkZg+WibacF+B0woQjK10eCOg6ftRjd0i/IraIOuV
i38W8CXGF5xxLrjBZM0yOV+OMnVVADVpn7RFDUAOuuvWZUTh0dYuNa2SQCYZDPl3
tCEJObCU0LhAZRDgOYofXk6mTqrbdepJWrb3GkEW9VuCghg/qX38qXqdtUM19tCq
kKYDXLxzqnoqtlhsWa/7CAEdgFbP9RYDU8ZxZzkA+3JGbzdto+HYQZJlhmQBNXiW
gVwx5Phr4jOWktDbahfZM/190yZ0bxYkHZFdGAvN9UVlT830r0ghJ3A9glMPEAD8
cqexGhpMX/nR/pNicLwL2NJCfrd9dNcwr9Brp6IBN+p/tvlLU9bUU/vm4gamA10a
5DMSaxjSjDqNnXW3KfFd5DqSrsEVrBYXnFKC9HaYqMvxaDqb92+kvtQDTSdeuP6G
tqItaDyVfDX+ga39waR2y0xMdF8OiIbW9IVtn6TBgNhSoL7cAcJznRUD863YVenI
W/FdFH7etLD9A1uixsipY5cOGf1oOjpXYTJl3oDAq5z6MgPo5oPG4Zr+ST3IUoez
KNz5HbYgGUzsDwruX+qVjcGsKW0jEVEBgKpS2WovxVEnYLJ+dvC1+sAj0CD4sej0
AMTwiCq1BNU5zg1DNC3hj5RHTwnN956xH4YJK58nwdQIxiJ+1EcfWBGpp4y56fiX
Pm9krKJQrBuD+O+a6JH6PkuzGoeCMmNudAwV3oTuYDX6/1uGKTKDwLK76fDauFYa
KnGklhfKyg/ieh9ItKzTO5ZX+jzd0e8dBcKhs9syFNbjrbqCyKOo7DMFrXu2tRw6
WIMoXK9mBxtVySo2m8BdNzgIMrA9thtti2gNSilMIN+HneX8ve1zOsC2+coz7Ri5
ZGyy6mQ7IyAM2W5yf7jBiaTmOZpwrk2o+y3nbgyFiS8rDoGlBgjLV0FD6N3yZfem
RWRJZrkCaJ1Bj4zD5oDDZQAZOO4AAqA7VDEl8fNCSiIV6JwZlmfUres7k+Ew4M7q
b3XJoEts1BH/SqNDyCkLr6OCo+MkXaJLgv/zn7iEYi1lVdqEIVoAZy/cw+Vs3w9p
TT4L9jKngqvbOdts3JQqud5Rek58EfdKYuP0Dl1z3mdYoOY+xGgDs4+v5/SkHTzy
gDsd5HVTgx4/nxVHjTY6nToGtaGb0l686dHRtkp0Fwv0hAhhCPM5VKVbzqNmdN89
b5WJP+lxo08/bxJJpcasi7nRp4hWKGqQKPULm12g9prQB4/HF8OSfR/M4iRrQj5N
FEVWK0E33VbuT/gsguG9F6VJ560JeNjYh5++h9hO4tLw1e9FOqTF+xmx2xIcwGCe
W+MBXbxD4ottObw1A83H0oWnuS1nH1f+bNT2gtmIcC+eMWVqV+xnkY0Af+NM/1fR
48AAv3DtyXP1tdp6ucqL3CsBORms6wfgM8vUMN5q8YK07nbky/DBa54k/tHJiNN8
acKJ+AJ+U00CXAPxdGuinS04Z6fvnZBF5DrGn2/sJUCHzMra8OcxcJCG3z8u3gJM
vNBLiUos0BTk0vVJ0yGbbTJtikF6YjjcCuzHnmzBV0tmQAK4lyC0FDi7m/0RA0mK
fRYjOnI/5YWt519Bp4PqntG+oW5uOIQSdXYO7WvBe33WPI5BiErtuHoS7nGhc9HI
VyOtPD157vHjQZferpLbha0iPHZcYhv0ao2LOdUe6Ag2hny/Ht9NElkvMOCbwb89
gOgWbSq58r4X7sbI+wBnnlt0M1Unn5UjVNJsfu3mbJAn/ADMcJD0jpf4Av4dIUU6
heYjV5+5/wm8fVaGolTvzVsjstRrw7R/OWxf6Pb9PCTEyKGCPApJF6QjB8CQUctb
98KmKUq5lB4maclr2bqx0gn+zWgeUczle4wIeBwnDjM7x5TYHBLRhzOW8/I4mdSl
3Yx4daSUTkW4xU5BpqmO05WerH1tVlMMZWqNxi8iYAkkicEjhris6MYhL2UncUlK
trRMJ8GR+etSnCkS+x0DIb5zU5YLBvnwil1xTpiarkVVQMcEoove8EDut4nSOo/O
drGUd2PBvL5m+1ch5ydPUoOnXLRpCOn1z+Z8jSAjNM8Fi8B3eSEKz3dd36V1x1SV
bDQrqOiFs86ixhrrWmXSVhcwjA0vrG9ByBcwSEEH8TXbKo9lk75k9PPmYb0H5N+3
3gnr2KLVmfY3Wv9wkpoLOJiVI3x6mpngIScROasssx8eo2mKvMwQ9RVHMyhfyRmj
OVt5cifoBgLRPSOJpFiCCGEet7THhFDXdGEeLSj5OcE9os72FffqDmkHngE3a1ZR
ZAN0KxSH/zH3FWJEhZZjYr6tYxCYFk/vXrMJqPmtCwI58CWqNrgUYPCLkyT5mlpn
LiOKa9JOVziwT/bW6TwqEmk4KCw3RIyWlVJlOR1vpPLotyl6ANEOGEZsVOgkF7Y9
qPvWqOFX/Mj1u4ixPhnjiG13pOVhmQvy1a97mQJmxlNzxjTh6pPCKc3SmugKLX67
NtcYTPGzfJ+AcvmA/q4mQosMP3QJSZE2xJMuZWFAD0SgKwUSEIybmy9zTPPq1OSe
G9NbqTyiHtPAFDLx3T/qCsWuW/nq1Gk4M0FfHiChERdoWDeIGk/OtrvN1EVIBVUV
UjSiatTsgT4VyU2HSkL0vPC3iZUgFSHKtWBVhLdP7RTEmn/WYQFdLFDcBe2XKcbl
zmRqHqG8hO9vKFS77doe2D7XAYkVml/96v6qq0Fs5KHFE73mU29BJ2dtKH5UXT4U
zE9yTzVWFbdWl45/2KwL9/lQx0oFHczVNzluGoAuOb0lATnkhPefFfjG/dYwpnID
atTi/ZUvjaXgcQVf5ZYcODPvhGhQmeNBCcHkr9rjORDnFufYNw2l+rbUq9Jkvor4
S9wx8zPB7l7++R8pAgo4/DP/iBJ0KIZ4cwgx9NdlrrxKRjvnoWW0TxQheHfuBkfW
GpaOWkwydFHvhVMDy/csjtey6AKAW4ZCb3mPPHyKH+LTr6fsV2lU68t9WdIHsQbh
4sWFQiAdyuw9M3PYbzwCpPWJcwNWdTXiaI2wqXd+jjjJx3L59gvKCi0FXm9VdoHh
Ap1E+NsYeFY7zwvqLtZAeWX81GNjdsI4b3rGI6zM41O/K1Z7WNXN6FaGaDhw9/gB
trCj8xvt8jqCcyeeN0KXRO021uDSYBomQ3OgOnMAcmtIW1vZ3/uAYt+rKZDGLn2G
sfNd0KfqnzI8EqRskolFLZTUBYlx4pp0Pa9xa+f1QBU4KbS0VN3Z2Qspw5vE8FQk
apr+hGFdaqjFkaJgPh5OY0k06G78c9yym9pN4Lg5o/fkp6ExGdGvh3zBYpjrMS1J
QdX25NPWqCFH8MABJkfPKTu9uKs9KvqqzAHCC9o31C8cVhENyDg61oq70epFHt5Z
TMR64UfxdT0KpsPRK/CqrmvHdD/pOL67BCvQRo93vOG4NzzLy+XmVbz0hDRGKqlO
gHwx0rgL8/za32K8TX9Xy9EMKTf1Y9bfrZSnhh3wg2XUje18I0LAtdwbYDQaJ2sS
CLCLN7dx0FLifOAjXN67gNug7w340Q/3rOapgFnnWVj7FhTwzUj2j4MECTZNwl2/
F1DkVTUe7bBXq+UMAdmYCJZ5WDHVy3RR6XixezghD15jLu4ZmBsjdwdtNPaVsJu8
nz7UsVQlvGlKWI+sVs008+LzBFF9gspQ0LRFxp+KNqzuPrq1hWKvl0Jzc2/DaVA8
CwpWvD/+MGUDy5vW2IfXwkD6UyUmupAVrcOpzdJEvO9vVEaaK3gOMM09/m2CdoZY
8OROip/TVjNbZ9/QXMABi4x/T71a6joaRYS5Yc/J1z0Y4FAHzAjyv1h1IPWcNrHB
GF/ND5sKcCBzWC1kQeVmbmffdlZvsXjJ9QTGjzO37klOVavGRWBmJGizAwdIhc0J
NXZokQB5kKnAhJd22MkS8/HiwIbOf8FNKuS9sG5eykwbvgrA/mfJWB47OOhqxERD
W1Nt6arGO2rmGI0o0gH9+euQinWgOgzLhWoie8sHZIChxW6l4FiK4i2diCe4hbcC
ZuEVGZqKIiljY/AQnU98SVglrhzBuxgB38EGbpUbc1GuHBUxVGOlT++JUYcEGcfr
sGGKGGiPxJ+BxaRgaenprNLzEt/Dl4A5YCo4gH5FM2kn09R34KXyf6dn7LjEzfuJ
NQ7hR6LX6SNadh9QkWyGEdJwehMzpxIjSPQhmMH2GwJZ2k//USDLwdtoS/W3+vPg
LbtLW7TrESSD3MRW2f6HoJvAQ0VhzyEtMh9Vde7r8OK90vN6L0iOKCPrHK4aQCuh
D5sNr3fWnvcs9YFgdP4wYF5tsg4cMj03p8N68WnmXMImgMlCwPareDT9/voHTQJZ
XlFsaaEUc7dI06maCkNEvV9oFh6t6zyIZ9x+B8YlX6WtQINOtetkbupLMkQ9k4T4
+cCqhOZwWm5DL0kSoYElrlDUiNVSziF2p+6MUVqvyn/AXnQG3nRFGquGj2OIcm2J
6DRPE/RiRjoImd2vHkyJ7cb6CgzwqJoY5MesuyDTtINgbUFckzOJyH6ezCbWPfdD
vOKxQBwa2oldmvmImhmimIO/2G/ArANQxMCCgx2YFINX4cETc7guWFTWKUTIb5vg
rVz08v00VQh3lLlk7+LyUOr511oMKrL4PUzBHPiRAjqC5IarGF6YbBCFVZW9FJGV
piXIVUW4dNJN+U5YQHv4+qh+TKEAn5SF9qtMLSmkpSHN7+cYMP3FgTFsz2Rpfa40
kekuBROBk7KC+heFrbTvCllpL5kFelXxegYLCyEAlLx7/oTAt3iYAx5dV2R1lUCl
r2HeaxpYDADvDBgAqsZCScpnVyE3Oj3jU+jn30PrUr+z+4xcZgf1wJMdVYRZU+TX
BPHeH+i83YIn6bhXtbAZ1+FEKYWokQnZWYIvXMI8Y61C2qJH6eixXJy44sgAto9K
4+A9/jY5GhOXEQCL0xW3mxEbTrpDL7ZtjFjubfKMYNYETzlV/CrbRwNE9YDegtYi
1Cb0OwOMHKxyToZW/qAZ3EvlXC4huxVQSIhsjse8qrMzUIAwhXomq/KfVRTmQaGX
IJxYUF9/wITKWTd7dwh8N/K/LMc7DkbPVEW6Vu2Y++R3kp4cClpVnehwag/m9Sim
woXhf2oaksT9s7kBYwYZ5X8oTMm/RGu+BmzYxK3EmF+jtdo0sbgqyDcRuPBU/pFL
9O4OafeVYmYXrUihise/BX2YHvFcS18uWXSSNgwHrk1w8hYJQTYOyNmA7eGsThcO
x9TatPQS48I3iWDWagKSYv9VLYNLAvzrgRGWjyRW0lzbQQRZE4O2om+4BoChNcYS
EY1B/sB/i76xaTnp4xpOO+JYiaEuidz+muzItz6qEA+cYQGwYF9O4fAO75UT0TpP
2mJXlrWvnyWl8BVuNybuIeWK97XyTqDm8IQr0ebiMmBasbFPIGZ4o+5BwxRHXtw5
XRmFhChfpcAOpZLpyyNpyqACR4hZfzgmeHidqrJ/QNdbTUIhI6fOmsqzx0QYeX8F
LgXO+0HCk+WBE/kwXpGs4nbROh/ZDMmrk6CkFhk1MylHzPQONYltpfF3PIC8Tw4W
VLNkqfq6r/NZ3f39pO8R1LzH5FaIO6hmU9g4Ze0xbvy+u661q9OkAPCDfbG9z7wh
dizXwSIjGVr0L81DJz5FPhWVGg4oxpQ6rU11jZ8Rb2Zi/8iH4wLWABrA8kD4+XtB
o7Rv8MQxsSP99k1kw+QlILNbWRCdaEpBZudKsBVt3YKNJ4oZEFKu0+KoFYvrfS/m
iaRc4iPMRgozvX3+laTu2fePslwDM6NCXMzCbDY2zXXXnsx1l++zKJ6kqFJlZQ5I
8wX1XsAbNCIQ32tDh+T3UrBZOXzI1FWNDAKcOvBrQ0PJEwdhTXaiYIh/H1pQRBFD
jHahx98V7CLEbh8EUV5WESLgXvHmseLQuDxpFehNurswbM+iMnLQ/WCoNj0MN1vb
NqQt677LnmQfc/PVFLKgWjF7QdUUNxynhvEej04Y4YoQ0HP5dbs9AKAXMeGXn3+O
A6bWIHUwdxRzRMhF8040ytszXvkV/aM5Ir59r8GjIlB3KuxGuW2Vto1SWLCgjzxq
IiGoCZn10iT1wz5aYuncVbF7KDACbHvLzuRnyIynuDPremCPzxs2/z+FuIJdryko
8XgK/+yE+IJuXdjBlm4ZAa+HvLX2QOmq1RWQ2xGVtwbuNmv7c3V5kQinRNE4pyO4
PztM+hqnPFWyYO9C/4FSUoT4pNFDRkVuNoP7/C0UIGsFuS9rIyWF23tSvuPHaHjD
+gjm0pvwjBw7OlyeIwlUZ68rBtQSP+0PyOO4y3h7ebmkfLfDCs6DAPp6y9mGtbAH
9M77TYKivfO+CyDnbOQCM/gxd2gphiF9khxFB9fxZA4LgY0E04gnSSTQrqkbSwt1
ts+UdGS4wHKpOLRKGRUa+ZNTrc6C+Mrjpzd9fBLXqtgLG5yCYIdqj8sDhDzn8UuG
RaDZ7Md1n0P0NJIboiI067zoW3+uGTJ+gSa09PvPU0Qz9QVozkvUDFLjRbs1pDxD
0OxnnsQJ9mOjvsyGq1kYjf3o0Z+0wVBL6GYwqQJR7PJm/63Tnq+mtYCFGPdKXXfv
8JGDf5ooyOZ9DJJi2U1XuQrIRhzTvH47jlxA4agIKMWJh72YNFYbIntCMr67EJ3z
80YRHq/Kfq444JaIGW8kRVTtq/rXTck8iOGwA027p6wwRqXynEYhkYBYGGHtmSxu
GdsiBkqgNqvyoQuFFfPWmrui9d4IMKtcX4DYtjyGJ4zCAsMPYnlQG+vS1BwRT24y
xd+jrdoY6iVpFh3SJq9mqhgE9TSEUk1TB5ve/1r/xV0r5M55vfM1TDRiVg1Rws9/
C9JvenNXbVSHWcyztlcpgtJ/LG4sazRLWr3qUM158ojiDTHuYhXIxbMZFCG8mqS5
5HFCOSf18kdl0UKbzEy7NU5h9bzau0mlAKy81KGUTTAYmvVcsWXWqOK251IaQ4mv
GFNjXK8mkQlQwknrn7GaBYQe/cO5p6tvLkb0Ct2dnA7mZLQPzyGvaREcvQLyUM/H
j9dyCM5R7pGpfO41juc+WxNKXbTIn1QsHYOiyJKF0kNbKdCqLmIPLxlXNK+Na8Hf
nVl3r+nrfg7EfG3RtqB7L83afL50UmpeCOZMnfqCoLt34Qda14JgAVhkSDpdu4o0
abXZvKxduuazeoIt+N+X4MMCDhFYwUcDTdOX1ROBNg/HFJb/LGIEish4qKLZRLLz
KQ2GoYEVHplRqWJJTC0HhoX+VBTwarzSr8vQ3CVpRr62R0rkzsx4XBgCp9ziDxQ3
jon2faeyvq0is8guCNqwKBL9iMt3zF/Zjms07V9MyHBYE80Ilig2AWbVNoSZwFOq
2J1KJsdGyP7HyHb5w/ygk9eivH//YtF9LQHmyvFSUXb9vZpJTYji8KXIMLxiMGqP
WQAB7QAA0OoN4vXExNhWSp415//2i1NQLA3PoFpofcRPtq4hIRtxs6QdqXG7QZAG
gnjBoqbPmk1CqjTZMzBhi868XCP1O2k/klSUEA0k1PmnDdQgUwZpeRRy3qVXOwAq
WVlmaJdzAPBfo+V1X4JOgsmPAOkXXZRGqHD2ZljDrVe5pZgVoHp0F4duv2LeQOJM
O37IruDgLQF+UFf+lqksuGNss391aLrU99dYkMk3PZsTDQjVTzzyS9zVgUH1rA2v
YhoWEEXub8LU0WIz1/WQNTHakLXwtdjIGQSgBNHnpb4mNyMsUmy7sC9ZGvBis3OS
t4fgXUaJsfIDYXRWulcz7yo94T+vtQ5ljIylrlw7HDZMcNRkrHfIxZ3t5Qz1GCP1
XX56pdZPki8gkkquP4NP/mbxk9E51EePaYeuF3HOlGeQsoyRXDNJSQHcUzBiOU+w
27IUwgmEOnLFMMQF2MdH7Z8luF2our1y/vAKQ4s/pWITtQcMy0lCrBezeLQsKctD
s60op5mUDoMp+bc53eZt0ClcYY5gvwfmS04LIqJg8FesSDJR+/4TOGIQyOyXZJZ5
UsjESXEgH2fSYLn+jUwLrKrxatDduDTJPxuC9aRhbIbjR8xlyapIr81eGqCct3ZH
iGVu4OlaWY1xGmttEEhy0oCC1m/rFQ83cuP3BNhgMXxCg7KhmUWzVvyFz/1uFHrW
IPX/td7uTarJp3x2EPauz04EQ3P4OfZvqV/xGSp5BeDbOUJ6D4P8xBSw0qkBVRDN
+yTAakOpNOtctgancZfiw7hhq2AjSVuCDlQ46GWZFJq+SmLL0/EUzga/6yNu2Qyz
4u1Wh2H9jG1Y//rH8bRD5eTi6lQLPeCH8fw6LkwEcq79Ccr6KzCQ6zi9LU4xGVnT
jM6s/yIWVV1nT7ZF1Ftmc/kwxUeZ+3bkNNUor6KNrCkU7+nYGcrsxfiF14nulUpm
pDRTbcpirChqQ/VYO1q490ddCQ/lDmLCXQaevU6yUiZRZiUx1nzm8qc5ixjXGUXq
lp1WOTKP4YulV+r10RqfLvLb+0/HqSxTdo4sFUKX6Hs8CQso9mJ9LMMY+4efWJ75
QVLZ0Z+8tJC6QPPPuYaFrtCwrRFC0P7uflh/SKAd/8TUBkKU8EQeQLbzqF1WqnpT
UQ4J36JjaVP4vbIqDHLkp51q3CKMATonyDnTZt2YKVqLt/rGLxsvF8qnuP20WVMz
fl1hzWy6cF6utC9LJko+FnfXyWOHm0UAN3qigR+nrRQ0H8dNMCWtngFQcvpAMaBR
OAzq5WXWHZ9Q6zaiQfuPeKw55dRS9+yIgFcE/cjopEqJtToOZrrRFSWOteDgrmx6
7ChkswVm4gmF3u7CZQYFnNOq10gz7mRe5KopwoARFvXRH2C77/n9PtZCNHmv54Kr
n2l/mj8TCI7vkrnvcxLWeF8brYbc4OEq8/YF0EhDQsUUy5bbV5y0aH2V10aBeKU7
AivigasDMqeqninjdzjTQU87/oUnGW3pJnELQXVN+RFSAuuULhIRtnYID52S+X8O
PS42dCobW0SDD977x4EdPpyxHIwVGwef7UAe/3vK3QIhkQq5tjRh6qmMgWyLPDke
wE4Kzgqu3X1hW7jGo2dvofbq8wzlC/ZzrQmW4miyJ1m8LIvQkRlfgDggdwa43jBE
5V6mwK97Z7CP8Z5EBjEb7oN6WtLTtZn5uegY8HcvDNS272iW6PX4IeKfi81Nv92z
cRK8LXPuSpD0Mjfe9OC+dVnmXwnqec19swAlgNTH6Ph8ZfkSJSyjzqYn5J9a/Q72
I6jezXRYi3nHIWps0x9xO07ekiTGgY9r/qjJLYzT8KUWWNm74ZSWXNOIkKkbGxFQ
7OLiEbmnleT1HuJgtaZbUTUMty0gi6Yox4OHjr9cwVK+vYjw547TKf63EQgghhNF
iW6GrXEhI80ZMYl9Tn22rTnl2Ph1xsGssYpcRu2tewJYoB6ySUwNfopU5kxIYuJz
/zhz6foHri4Pa7UeIyLS8Ej0+yDWqldTiySCjY27r5AqHq+RHx57w2nvneRqunEl
a6EbbFMAwF5n6qJ1uHoRYTC3gFvx87lvxBFhW4xMJdD+JAVVHQ+kYg34zgclu5cV
sqV6io4ChutsaSdMcNYRES/l0QEMqV5DbJOZlRtYNdIPQpvHKQEZndNS3Iyx4cD6
cXA7swii3nFpx2/hUK03ZOG9gKbEA/qjS+BvJ9C32QJWZXz0q9yy84ZGPWW2+PLZ
j0JKjJpMM9Xo/0b+WM7naE/9XZ0xolUnPqpCxJlSl4RKbLmgPuehG6ATETXiEh80
U3tUd2bdfbr3wW62VbhaPi54N9KrhUjyJaSlLy3qzrAI76FF6lBbQ+gOqiG+5htX
kpqNXIfvUrf7N40GIibrmdQkv6pgG6L0FE7z6JfO+3p4x/ev+iotYe/O5gu/jCVz
M1h8tOWodqwa70vYk/mW3M+o9+BcyG18IXfLVAtkLKZxPmcxlhRzaIONNZknszvR
9SqMrWXlBd0vqNpolJlHP7lkARa+zh5QBDU36YCe0xuH3RuUgqZ8Ggb9A7C/v4KS
p7HXyz0iTlr+Yz1VpMlTQnZdcwt256Zfy1+Kik5O9QGcKZp3zN+9dTIps36bdsdg
RO8RWc74d7gWwO5+2oCHK/7Qd0YLRu/frbgwLu0LsQYnM7eFDrFXHxoLkBh1V/gd
WLfl8s32hmR0a0qrKh3KC12La7+2z2hezAGaPQq1ujtmKNqOZMHC2HwankKYUqT3
y6GbLLUbVg4YecWRomLVWD67ayliowvOcNEfgnAYoShRH/nYHNbllC432+CVU4VK
EeV19Jj4ssF1sA/9s8WUK6wuV6+6HxGNgkkBmwZKJoUdGoncSyl9pP+j6OUG1lox
tP/az1kvm7MA3hB0snw3nlLv/ozvXkiMZJ3vdg4KWd87xUCb8XlRlCOFqqWG0Bgz
WMi2JurMMxqUNzycwExG/jdTN83IZqDj/5q5sMWdlSUnpnZinFsskPdkvoJfDgu6
EMbtfKYreF99gD0r3ORAWy/4NCl5r1BXnUaRvsncPs4oiUtxZ1RXlnPpHmgjb7oj
GFjf3mqhaj6i5oHouHDeWpv+ZX4Noak3mK8fZq+6MabojZ9O8/XYSw5KJH3fPgBq
+oLkH3V2XUNobzvznJ13xImO97dhEOknKuC+uiqKOnI6kqspK+aaCcD3a1fILFDJ
XKRE/FxnfCdk/yCnYJgPRxUv0rqOHHtDNNoMkWLB0Ug9frIO8zLFZfXaAXoTKPho
4uWDMlV9dVAAixxfDZ0iVo4Vjv8vGn1PlClBMtbVtxy4GO6YaITgZgtGpbbTHLcZ
yeIUlWABn48kynUrVb5uwYCse8gZopogN+IOr7jwO7bx7bCuXgoCEorBrhYhV/Ht
PPzufpsa/stdp5CMM3jKVz9scYmwznYrrsVVEOimmiHtzsm+jRjK05nIQixxPfh7
dWMbSNAZG643xPsmorWKLN9Ssiq7bJ6wthDqdtifFEsxdqsIDZO6EhgpV57cET3b
KbQ9CoG30xj1J4e2nD0I5v5fWb1/FOGxdshCjwPCeyCXKhR5OcpLfqrnYByIJwoS
zljt93jrgwv+hL+H1fB3pWztuziNHng/KnaX/oHjFqKTK3K9/yRhMfU9cxUPLxNB
Afn2qz4rCGMsWJ6uw6L2W+/ylW39CpxQIkuJcjGCxy648W2jRWx50znTdPdnjnWX
dWyr3rVOVWWeIS442hCiCTK6LuSyaOk7jZOIr5bm6ULoegsvWtI6DLrnGQei9dLq
w5Qub7PImePwfQHqXULFJGMP7zbhGXDH+cRoNMJGmO8/rt0tMvUcpTtdfnCH5jEn
r9DB23dCFEMozRMqWOEBhKKJ0lUSQ2U+U44h8w2FJ/p8A4xv5tJ6nQknVggytE0v
PqMtBvLq9SdcQrvNzb7sZ+RXLWPk+06b14n5wXQ5ZVvFZ4PL9JvZltvL1TqUT8ld
gAeJ628BnA0TElWKho1+8xvk1sFcjojoqyhFTyPSVLEPmU4ctWF1fzz2H/APCPO/
qZG6yv4qseEO+YzNbBquOBnMdZi/iqKl1ZLtJk13fPX9WDiErseu0a+4+oBTmtZ4
hi9/+tsC1p2jqUvvwjta3Ti4RnFayFRqlA/0KJohzP9vIixzRSGIQAp9PpfeBG/f
OBi3JJfRc0OLkMx/+FIoKC1jhiF247wMN2wc5BK0rhXP/li5ucWDrN1W5MnM038y
w8z/JLlxx5cBOrMbt0pktVcxJDyRSJsVE8G0lEf+kOO+RI8eaEM8gGBoj/dqOQvE
gWJe9WXjLogC4Geu6GsioAIE4v7sDvvK9LCeEsheGwOjAMUdlGMMFcQ+BpxOWXX2
apfLdNU9kXQyk8Wn6yQ6xdHhYvPasL7ayTdi6d9iXOV8MFIrb7yEJTfGlMUY/KJM
UdUMvU/6wD47nPC59JkZkNbnubM7x1/rpq48XgZT10o44rsQnDhN3AgKHxGv3zni
HgP9kHPUW88ysKJvjgfscR9dA30EXcVcIuEhJ90m5H/siDRnciwOUK2Ty7fDnvgF
6zHqzmb46GSxxHBeQsBysnJ5EUG/a7+heQf/mScWlgZeF+jh0AmkSg5ptMmLumfA
6yVNPQ8Ziq0+d9B4EZHheMSFIzSqBmDzLmQkeCYpIFNrSjHjV1DP9u2xJ0W2FAps
Hg6tlhgex4Q0MJwwuvadHtWBemMuOs3bCGukv3SJXSVhedjjDBimKyyifyg8ZoBG
ILP11wCrixBAlwL6L5UD3IJ929eQ7ZsUsfWu+CS6UAfbRkUIn6CSuWrgnHClfSME
h3VLqmB4wLOGL9fy5AZS2sZ1PMYPZ5VrhAT8oKYxqV4vMXItWdPd6yi34bLCXE6T
+YmykjmM8wiEIC5SKcDvg5460GZ7cN/gOW1UMD5yHfBC3E7YltVYjqHl8G1dpI30
oUvSsqkSNbDOUGjFH/tDUWrCxSll8EZGrXacLf6YQi7XJffJPp1WydzP59apXq98
w+bEf1z5JpaV+rbh5x95A9Py09uL4UNu8LQ11LuRDVhiy7GGAMfFAF73Mm3z+BPX
slJPblEe+apv8AuFu9U4gP5AZ8aNvxhcP7sLBtNVCwggwRk22OaIgiNlEJ9z3TTU
R2TFYs+kR/pxhV0BgQiJkd0pGsEEAPj25BGl1PzMQyenFTca58qp0WtWx9YQGKe3
Ho95jBXLNoaWaoq4WK9YOy4FOMggDqB/+hpDWqW3VQx3ZWV/2wkXUE4DC9VGtPUd
vfPWkgD5ci9Mk8DTsJCCjjqT1ocIe++rSb6OziAMUNw6Rj9ryQO3mLzPj0afqiV5
FQ+VZWGNXRDQ4rK/rffmiEwgLdGAqwCDb5ZmYJTXLilNJ40FZmiTo90hELx9aM0+
7hNSwpKlOGCPjz0q8dF77v89T92wl/lSUfwiFy5JZHt2cf4nvGyCOFtYNVN23P5R
+0scnvesQoct3y9AVPMzRjcMvQaxDVgdXtj31vFm0XVNrl5GN2axHOKeypH6V9cP
kBVhkZ6QPLMS3jlQqYEkk+331uTx9mRduOq+0LyR4seZo/3N0XyPw+020XjqcvAr
JHzW1YrxUE53SrtmhkC2Ogw5WQZPWHlRkjJeKTSvkHM1ZAc+rH8Ek6mbbVXaAvyr
WTLs1xfXBpnGBD0cf3/tsxjeLa13Ssc1slk6RLwBdzaSBF5k9k0+c+iaI3I1JV44
J66SEFxzBnnI51wIY3TeIGjCZD5sq21P0bcvfMnBlQh5on3f5cMrwePU+618KPlI
D2RAD5yy0H/z47sd2SF8uIW6o60hCMT/+xXqTgAVth4wgfDqB0Nosv7+2sW2fxZi
xoEqnzmKUq8jBavEBSROHlkGavFFcFc8W7jVqt8sceSQKnNzZMKSpfptEezYF2S/
NgHzyAEqtCRmAoLGUf9M+3HSqB8E+RnivC3ZCFDMyJ63O58O5pe6wrhy4WAvDdz2
7V0E+AA3MI/aznLGeYOYu2o18b6UIAucaNDtDAsqNJw=
`pragma protect end_protected
